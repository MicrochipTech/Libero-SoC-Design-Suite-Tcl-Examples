// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAO0IlI
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAI0IlI
,
CAXI4DMAOIOOI
,
CAXI4DMAO1IOI
,
CAXI4DMAl0IlI
,
CAXI4DMAO1IlI
,
CAXI4DMAI1IlI
,
CAXI4DMAII0OI
,
intDscrptrNum
,
CAXI4DMAl1IlI
,
CAXI4DMAOOllI
,
CAXI4DMAIOllI
,
CAXI4DMAlI0OI
,
CAXI4DMAlOllI
,
CAXI4DMAOIllI
,
CAXI4DMAIIllI
,
CAXI4DMAlIllI
,
CAXI4DMAOlllI
,
waitDscrptr
,
waitStrDscrptr
,
CAXI4DMAIlllI
,
CAXI4DMAllllI
,
CAXI4DMAO0llI
,
CAXI4DMAI0llI
,
CAXI4DMAl0llI
,
CAXI4DMAlll1
)
;
parameter
AXI4_STREAM_IF
=
0
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl0OI
=
23
;
parameter
NUM_PRI_LVLS
=
6
;
parameter
CAXI4DMAl1OI
=
133
;
parameter
CAXI4DMAO1llI
=
(
CAXI4DMAl1OI
+
32
+
1
)
;
`include "../../../coreaxi4dmacontroller_arbiter_parameters.v"
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAI0IlI
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOIOOI
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
input
CAXI4DMAl0IlI
;
input
CAXI4DMAO1IlI
;
input
CAXI4DMAI1IlI
;
input
CAXI4DMAII0OI
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
intDscrptrNum
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl1IlI
;
input
[
31
:
0
]
CAXI4DMAOOllI
;
input
[
31
:
0
]
CAXI4DMAIOllI
;
input
[
31
:
0
]
CAXI4DMAlI0OI
;
input
CAXI4DMAlOllI
;
input
CAXI4DMAOIllI
;
input
CAXI4DMAIIllI
;
input
CAXI4DMAlIllI
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOlllI
;
input
[
NUM_INT_BDS
-
1
:
0
]
waitDscrptr
;
input
waitStrDscrptr
;
output
CAXI4DMAIlllI
;
output
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAllllI
;
output
CAXI4DMAO0llI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0llI
;
output
reg
[
CAXI4DMAO1llI
-
1
:
0
]
CAXI4DMAl0llI
;
output
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAlll1
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAI1llI
;
wire
[
NUM_INT_BDS
-
1
:
0
]
reqValid
;
integer
CAXI4DMAl1llI
;
wire
[
NO_OF_ACTIVE_FIXED_PRIORITY_LEVELS
-
1
:
0
]
CAXI4DMAOO0lI
;
reg
CAXI4DMAIO0lI
;
reg
CAXI4DMAlO0lI
;
reg
[
2
:
0
]
CAXI4DMAl10OI
;
reg
[
2
:
0
]
CAXI4DMAOO1OI
;
reg
CAXI4DMAOI0lI
;
wire
CAXI4DMAII0lI
;
wire
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAlI0lI
;
wire
CAXI4DMAOl0lI
;
wire
[
NO_OF_PRI_0_REQS
-
1
:
0
]
grant_Pri0RRA
;
wire
[
NO_OF_PRI_1_REQS
-
1
:
0
]
grant_Pri1RRA
;
wire
[
NO_OF_PRI_2_REQS
-
1
:
0
]
grant_Pri2RRA
;
wire
[
NO_OF_PRI_3_REQS
-
1
:
0
]
grant_Pri3RRA
;
wire
[
NO_OF_PRI_4_REQS
-
1
:
0
]
grant_Pri4RRA
;
wire
[
NO_OF_PRI_5_REQS
-
1
:
0
]
grant_Pri5RRA
;
wire
[
NO_OF_PRI_6_REQS
-
1
:
0
]
grant_Pri6RRA
;
wire
[
NO_OF_PRI_7_REQS
-
1
:
0
]
grant_Pri7RRA
;
wire
[
CAXI4DMAO1llI
-
1
:
0
]
CAXI4DMAIl0lI
;
wire
[
NO_OF_ACTIVE_FIXED_PRIORITY_LEVELS
-
1
:
0
]
CAXI4DMAll0lI
;
wire
CAXI4DMAO00lI
;
wire
strDscrptrValid_StrDscrptrCache
;
reg
[
1
:
0
]
CAXI4DMAO1OOI
;
reg
[
55
:
0
]
CAXI4DMAI00lI
[
1
:
0
]
;
reg
[
33
:
0
]
CAXI4DMAl00lI
[
1
:
0
]
;
reg
CAXI4DMAO10lI
;
reg
CAXI4DMAI10lI
;
wire
[
CAXI4DMAO1llI
-
1
:
0
]
CAXI4DMAl10lI
;
reg
[
1
:
0
]
CAXI4DMAOO1lI
;
`include "../../../coreaxi4dmacontroller_arbiter_mapping.v"
localparam
[
2
:
0
]
CAXI4DMAIO1lI
=
3
'b
010
;
localparam
[
2
:
0
]
CAXI4DMAlO1lI
=
3
'b
100
;
localparam
[
2
:
0
]
CAXI4DMAOI1lI
=
3
'b
000
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1llI
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
end
else
if
(
CAXI4DMAl0IlI
)
begin
for
(
CAXI4DMAl1llI
=
0
;
CAXI4DMAl1llI
<=
NUM_INT_BDS
-
1
;
CAXI4DMAl1llI
=
CAXI4DMAl1llI
+
1
)
begin
if
(
intDscrptrNum
==
CAXI4DMAl1llI
)
begin
CAXI4DMAI1llI
[
CAXI4DMAl1llI
]
<=
1
'b
1
;
end
end
if
(
CAXI4DMAIO0lI
)
begin
CAXI4DMAI1llI
[
CAXI4DMAI0llI
]
<=
1
'b
0
;
end
if
(
CAXI4DMAlIllI
)
begin
CAXI4DMAI1llI
[
CAXI4DMAOlllI
]
<=
1
'b
0
;
end
end
else
if
(
CAXI4DMAIO0lI
|
CAXI4DMAlIllI
)
begin
if
(
CAXI4DMAIO0lI
)
begin
CAXI4DMAI1llI
[
CAXI4DMAI0llI
]
<=
1
'b
0
;
end
if
(
CAXI4DMAlIllI
)
begin
CAXI4DMAI1llI
[
CAXI4DMAOlllI
]
<=
1
'b
0
;
end
end
end
assign
reqValid
[
NUM_INT_BDS
-
1
:
0
]
=
CAXI4DMAI1llI
[
NUM_INT_BDS
-
1
:
0
]
&
(
(
CAXI4DMAI0IlI
[
NUM_INT_BDS
-
1
:
0
]
)
|
(
CAXI4DMAlI0lI
)
)
;
CAXI4DMAII1lI
#
(
.CAXI4DMAlI1lI
(
NUM_INT_BDS
)
,
.CAXI4DMAOl1lI
(
CAXI4DMAOIO1
)
,
.CAXI4DMAIl1lI
(
NO_OF_ACTIVE_FIXED_PRIORITY_LEVELS
)
)
CAXI4DMAll1lI
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqFPA
)
,
.CAXI4DMAlO0lI
(
CAXI4DMAlO0lI
)
,
.CAXI4DMAIO0lI
(
CAXI4DMAlOllI
|
CAXI4DMAlIllI
)
,
.CAXI4DMAO00lI
(
CAXI4DMAO00lI
)
,
.CAXI4DMAI01lI
(
intDscrptrNum_Pri0RRA
)
,
.CAXI4DMAl01lI
(
intDscrptrNum_Pri1RRA
)
,
.CAXI4DMAO11lI
(
intDscrptrNum_Pri2RRA
)
,
.CAXI4DMAI11lI
(
intDscrptrNum_Pri3RRA
)
,
.CAXI4DMAl11lI
(
intDscrptrNum_Pri4RRA
)
,
.CAXI4DMAOOO0I
(
intDscrptrNum_Pri5RRA
)
,
.CAXI4DMAIOO0I
(
intDscrptrNum_Pri6RRA
)
,
.CAXI4DMAlOO0I
(
intDscrptrNum_Pri7RRA
)
,
.CAXI4DMAOO0lI
(
CAXI4DMAOO0lI
)
,
.CAXI4DMAOIO0I
(
CAXI4DMAIlllI
)
,
.strDscrptr
(
CAXI4DMAO0llI
)
,
.intDscrptrNum
(
CAXI4DMAI0llI
)
,
.CAXI4DMAllllI
(
CAXI4DMAll0lI
)
)
;
assign
CAXI4DMAllllI
=
(
NO_OF_ACTIVE_FIXED_PRIORITY_LEVELS
==
8
)
?
CAXI4DMAll0lI
:
{
{
(
NUM_PRI_LVLS
-
NO_OF_ACTIVE_FIXED_PRIORITY_LEVELS
)
{
1
'b
0
}
}
,
CAXI4DMAll0lI
}
;
assign
CAXI4DMAO00lI
=
(
(
AXI4_STREAM_IF
==
1
)
&&
(
grant_Pri0RRA
[
0
]
==
1
'b
1
)
)
?
1
'b
1
:
1
'b
0
;
generate
if
(
NO_OF_PRI_0_REQS
==
1
)
begin
assign
grant_Pri0RRA
=
reqPri0
;
end
else
if
(
NO_OF_PRI_0_REQS
>
1
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_0_REQS
)
)
CAXI4DMAlIO0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri0
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
0
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri0RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
>=
2
)
&&
(
NO_OF_PRI_1_REQS
==
1
)
)
begin
assign
grant_Pri1RRA
=
reqPri1
;
end
else
if
(
(
NUM_PRI_LVLS
>=
2
)
&&
(
NO_OF_PRI_1_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_1_REQS
)
)
CAXI4DMAllO0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri1
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
1
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri1RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
>=
3
)
&&
(
NO_OF_PRI_2_REQS
==
1
)
)
begin
:
CAXI4DMAO0O0I
assign
grant_Pri2RRA
=
reqPri2
;
end
else
if
(
(
NUM_PRI_LVLS
>=
3
)
&&
(
NO_OF_PRI_2_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_2_REQS
)
)
CAXI4DMAI0O0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri2
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
2
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri2RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
>=
4
)
&&
(
NO_OF_PRI_3_REQS
==
1
)
)
begin
assign
grant_Pri3RRA
=
reqPri3
;
end
else
if
(
(
NUM_PRI_LVLS
>=
4
)
&&
(
NO_OF_PRI_3_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_3_REQS
)
)
CAXI4DMAl0O0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri3
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
3
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri3RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
>=
5
)
&&
(
NO_OF_PRI_4_REQS
==
1
)
)
begin
assign
grant_Pri4RRA
=
reqPri4
;
end
else
if
(
(
NUM_PRI_LVLS
>=
5
)
&&
(
NO_OF_PRI_4_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_4_REQS
)
)
CAXI4DMAO1O0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri4
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
4
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri4RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
>=
6
)
&&
(
NO_OF_PRI_5_REQS
==
1
)
)
begin
assign
grant_Pri5RRA
=
reqPri5
;
end
else
if
(
(
NUM_PRI_LVLS
>=
6
)
&&
(
NO_OF_PRI_5_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_5_REQS
)
)
CAXI4DMAI1O0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri5
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
5
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri5RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
>=
7
)
&&
(
NO_OF_PRI_6_REQS
==
1
)
)
begin
assign
grant_Pri6RRA
=
reqPri6
;
end
else
if
(
(
NUM_PRI_LVLS
>=
7
)
&&
(
NO_OF_PRI_6_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_6_REQS
)
)
CAXI4DMAl1O0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri6
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
6
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri6RRA
)
)
;
end
endgenerate
generate
if
(
(
NUM_PRI_LVLS
==
8
)
&&
(
NO_OF_PRI_7_REQS
==
1
)
)
begin
assign
grant_Pri7RRA
=
reqPri7
;
end
else
if
(
(
NUM_PRI_LVLS
==
8
)
&&
(
NO_OF_PRI_7_REQS
>
1
)
)
begin
CAXI4DMAIIO0I
#
(
.CAXI4DMAIl1lI
(
NO_OF_PRI_7_REQS
)
)
CAXI4DMAOOI0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
reqPri7
)
,
.CAXI4DMAOlO0I
(
CAXI4DMAOO0lI
[
7
]
)
,
.CAXI4DMAIlO0I
(
grant_Pri7RRA
)
)
;
end
endgenerate
assign
CAXI4DMAII0lI
=
(
!
CAXI4DMAl0IlI
&
CAXI4DMAOI0lI
)
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAIO1lI
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAIO0lI
<=
1
'b
0
;
CAXI4DMAlO0lI
<=
1
'b
0
;
CAXI4DMAOI0lI
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAIO1lI
:
begin
if
(
CAXI4DMAlOllI
)
begin
CAXI4DMAOI0lI
<=
1
'b
1
;
if
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
begin
if
(
CAXI4DMAII0lI
)
begin
CAXI4DMAIO0lI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO1lI
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOI1lI
;
end
end
else
begin
if
(
CAXI4DMAII0lI
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAlO1lI
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOI1lI
;
end
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIO1lI
;
end
end
CAXI4DMAOI1lI
:
begin
CAXI4DMAOI0lI
<=
1
'b
1
;
if
(
CAXI4DMAII0lI
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAlO1lI
;
if
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
begin
CAXI4DMAIO0lI
<=
1
'b
1
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOI1lI
;
end
end
CAXI4DMAlO1lI
:
begin
CAXI4DMAlO0lI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO1lI
;
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIO1lI
;
end
endcase
end
assign
CAXI4DMAOl0lI
=
(
CAXI4DMAOI0lI
)
?
CAXI4DMAIIllI
:
CAXI4DMAI1IlI
;
CAXI4DMAIOI0I
#
(
.CAXI4DMAlI1lI
(
NUM_INT_BDS
)
,
.CAXI4DMAOl1lI
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAl1OI
(
CAXI4DMAl1OI
)
,
.CAXI4DMAO1llI
(
CAXI4DMAO1llI
)
)
CAXI4DMAlOI0I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAl0IlI
(
CAXI4DMAl0IlI
)
,
.CAXI4DMAO1IlI
(
CAXI4DMAO1IlI
)
,
.CAXI4DMAOII0I
(
intDscrptrNum
)
,
.CAXI4DMAIII0I
(
CAXI4DMAII0OI
)
,
.CAXI4DMAlII0I
(
CAXI4DMAI0llI
)
,
.CAXI4DMAOI0lI
(
CAXI4DMAOI0lI
)
,
.CAXI4DMAOIllI
(
CAXI4DMAOIllI
)
,
.CAXI4DMAl1IlI
(
CAXI4DMAl1IlI
)
,
.CAXI4DMAOOllI
(
CAXI4DMAOOllI
)
,
.CAXI4DMAIOllI
(
CAXI4DMAIOllI
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAlI0OI
)
,
.CAXI4DMAO1IOI
(
CAXI4DMAO1IOI
)
,
.CAXI4DMAOlI0I
(
CAXI4DMAI0llI
)
,
.CAXI4DMAIIllI
(
CAXI4DMAOl0lI
)
,
.CAXI4DMAIlI0I
(
CAXI4DMAIl0lI
)
,
.CAXI4DMAlI0lI
(
CAXI4DMAlI0lI
)
,
.CAXI4DMAlll1
(
CAXI4DMAlll1
)
)
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO1OOI
<=
2
'b
0
;
end
else
begin
if
(
CAXI4DMAl0IlI
&
CAXI4DMAO1IlI
)
begin
CAXI4DMAO1OOI
[
CAXI4DMAO10lI
]
<=
1
'b
1
;
CAXI4DMAO1OOI
[
~
CAXI4DMAO10lI
]
<=
CAXI4DMAO1OOI
[
~
CAXI4DMAO10lI
]
;
end
else
if
(
(
CAXI4DMAOIllI
)
&&
(
CAXI4DMAOI0lI
==
1
'b
1
)
&&
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
)
begin
CAXI4DMAO1OOI
[
CAXI4DMAI10lI
]
<=
1
'b
0
;
CAXI4DMAO1OOI
[
~
CAXI4DMAI10lI
]
<=
CAXI4DMAO1OOI
[
~
CAXI4DMAI10lI
]
;
end
end
end
assign
strDscrptrValid_StrDscrptrCache
=
CAXI4DMAO1OOI
[
CAXI4DMAI10lI
]
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO10lI
<=
1
'b
0
;
end
else
begin
if
(
CAXI4DMAl0IlI
&
CAXI4DMAO1IlI
)
begin
CAXI4DMAO10lI
<=
~
CAXI4DMAO10lI
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI10lI
<=
1
'b
0
;
end
else
begin
if
(
(
CAXI4DMAOIllI
)
&&
(
CAXI4DMAOI0lI
==
1
'b
1
)
&&
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
)
begin
CAXI4DMAI10lI
<=
~
CAXI4DMAI10lI
;
end
end
end
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAl0IlI
&
CAXI4DMAO1IlI
)
begin
CAXI4DMAI00lI
[
CAXI4DMAO10lI
]
<=
CAXI4DMAO1IOI
[
57
:
2
]
;
end
else
if
(
CAXI4DMAOI0lI
&
CAXI4DMAOIllI
)
begin
CAXI4DMAI00lI
[
CAXI4DMAI10lI
]
<=
{
CAXI4DMAIOllI
,
CAXI4DMAl1IlI
}
;
end
end
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAl0IlI
&
CAXI4DMAO1IlI
)
begin
CAXI4DMAl00lI
[
CAXI4DMAO10lI
]
<=
{
CAXI4DMAlI0OI
,
CAXI4DMAO1IOI
[
1
:
0
]
}
;
end
end
assign
CAXI4DMAl10lI
=
{
1
'b
0
,
CAXI4DMAl00lI
[
CAXI4DMAI10lI
]
[
33
:
2
]
,
{
32
{
1
'b
0
}
}
,
{
CAXI4DMAI00lI
[
CAXI4DMAI10lI
]
[
55
:
24
]
,
{
32
{
1
'b
0
}
}
,
CAXI4DMAI00lI
[
CAXI4DMAI10lI
]
[
23
:
0
]
}
,
CAXI4DMAOO1lI
[
CAXI4DMAI10lI
]
,
{
{
9
{
1
'b
0
}
}
,
CAXI4DMAl00lI
[
CAXI4DMAI10lI
]
[
1
:
0
]
,
{
2
{
1
'b
0
}
}
}
}
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
CAXI4DMAOO1lI
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
else
if
(
CAXI4DMAl0IlI
&
CAXI4DMAO1IlI
&
CAXI4DMAII0OI
)
CAXI4DMAOO1lI
[
CAXI4DMAO10lI
]
<=
CAXI4DMAI1IlI
;
else
if
(
CAXI4DMAOI0lI
&&
CAXI4DMAOIllI
&&
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
)
CAXI4DMAOO1lI
[
CAXI4DMAI10lI
]
<=
1
'b
0
;
else
if
(
CAXI4DMAOI0lI
&
CAXI4DMAOIllI
&
CAXI4DMAIIllI
)
CAXI4DMAOO1lI
[
CAXI4DMAI10lI
]
<=
1
'b
1
;
end
always
@
(
*
)
begin
if
(
CAXI4DMAO0llI
)
begin
CAXI4DMAl0llI
=
CAXI4DMAl10lI
;
end
else
if
(
CAXI4DMAlI0lI
[
CAXI4DMAI0llI
]
)
begin
CAXI4DMAl0llI
=
CAXI4DMAIl0lI
;
end
else
begin
CAXI4DMAl0llI
=
{
CAXI4DMAIl0lI
[
CAXI4DMAO1llI
-
1
:
11
]
,
CAXI4DMAOIOOI
[
CAXI4DMAI0llI
]
,
CAXI4DMAIl0lI
[
9
:
0
]
}
;
end
end
endmodule
