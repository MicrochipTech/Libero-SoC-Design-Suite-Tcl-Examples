// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAllOIl
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAOOOIl
,
CAXI4DMAllllI
,
CAXI4DMAII0OI
,
CAXI4DMAlI0OI
,
CAXI4DMAIOOIl
,
CAXI4DMAlOOIl
,
CAXI4DMAIIOIl
,
CAXI4DMAOIOIl
,
CAXI4DMAlIOIl
,
CAXI4DMAI0OIl
,
CAXI4DMAlII1I
,
CAXI4DMAOlI1I
,
CAXI4DMAl0OIl
,
CAXI4DMAO1OIl
,
CAXI4DMAl011
,
CAXI4DMAI1OIl
,
CAXI4DMAl1OIl
,
CAXI4DMAOlIOl
,
CAXI4DMAl10Ol
,
CAXI4DMAO1O1I
,
CAXI4DMAOIl0I
,
CAXI4DMAOOIIl
,
CAXI4DMAIllOI
,
CAXI4DMAII
,
CAXI4DMAOl
,
CAXI4DMAlI
,
CAXI4DMAll
,
CAXI4DMAO101I
,
CAXI4DMAO0
,
CAXI4DMAlOlOl
,
CAXI4DMAIIllI
,
CAXI4DMAO1OOl
,
CAXI4DMAO10Ol
)
;
parameter
CAXI4DMAl0OI
=
23
;
parameter
CAXI4DMAO1OI
=
12
;
parameter
NUM_PRI_LVLS
=
1
;
parameter
CAXI4DMAI1OI
=
8
;
parameter
PRI_0_NUM_OF_BEATS
=
255
;
parameter
PRI_1_NUM_OF_BEATS
=
127
;
parameter
PRI_2_NUM_OF_BEATS
=
63
;
parameter
PRI_3_NUM_OF_BEATS
=
31
;
parameter
PRI_4_NUM_OF_BEATS
=
15
;
parameter
PRI_5_NUM_OF_BEATS
=
7
;
parameter
PRI_6_NUM_OF_BEATS
=
3
;
parameter
PRI_7_NUM_OF_BEATS
=
0
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAOOOIl
;
input
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAllllI
;
input
CAXI4DMAII0OI
;
input
[
31
:
0
]
CAXI4DMAlI0OI
;
input
[
1
:
0
]
CAXI4DMAIOOIl
;
input
[
2
:
0
]
CAXI4DMAlOOIl
;
input
[
31
:
0
]
CAXI4DMAIIOIl
;
input
[
2
:
0
]
CAXI4DMAOIOIl
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAlIOIl
;
input
CAXI4DMAI0OIl
;
input
CAXI4DMAlII1I
;
input
CAXI4DMAOlI1I
;
input
CAXI4DMAl0OIl
;
input
CAXI4DMAO1OIl
;
input
CAXI4DMAl011
;
input
CAXI4DMAI1OIl
;
input
CAXI4DMAl1OIl
;
input
CAXI4DMAOlIOl
;
input
CAXI4DMAl10Ol
;
output
CAXI4DMAO1O1I
;
output
[
31
:
0
]
CAXI4DMAOIl0I
;
output
CAXI4DMAOOIIl
;
output
CAXI4DMAIllOI
;
output
CAXI4DMAII
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOl
;
output
[
1
:
0
]
CAXI4DMAlI
;
output
[
2
:
0
]
CAXI4DMAll
;
output
[
31
:
0
]
CAXI4DMAO101I
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAO0
;
output
CAXI4DMAlOlOl
;
output
CAXI4DMAIIllI
;
output
CAXI4DMAO1OOl
;
output
CAXI4DMAO10Ol
;
reg
[
7
:
0
]
CAXI4DMAl10OI
;
reg
[
7
:
0
]
CAXI4DMAOO1OI
;
reg
CAXI4DMAOOl0l
;
reg
CAXI4DMAIOl0l
;
reg
CAXI4DMAII0ll
;
reg
CAXI4DMAlI0ll
;
reg
CAXI4DMAlOl0l
;
reg
CAXI4DMAOIl0l
;
reg
[
31
:
0
]
CAXI4DMAIIl0l
;
reg
[
31
:
0
]
CAXI4DMAlIl0l
;
reg
CAXI4DMAOll0l
;
reg
CAXI4DMAIll0l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl11I
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOOOl
;
reg
[
31
:
0
]
CAXI4DMAlll0l
;
reg
[
31
:
0
]
CAXI4DMAO0l0l
;
reg
[
1
:
0
]
CAXI4DMAI0l0l
;
reg
[
1
:
0
]
CAXI4DMAl0l0l
;
reg
[
2
:
0
]
CAXI4DMAO1l0l
;
reg
[
2
:
0
]
CAXI4DMAI1l0l
;
reg
CAXI4DMAl1l0l
;
reg
CAXI4DMAOO00l
;
reg
CAXI4DMAIO00l
;
reg
CAXI4DMAlO00l
;
reg
CAXI4DMAOI00l
;
reg
CAXI4DMAII00l
;
reg
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAlI00l
;
reg
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAOl00l
;
reg
CAXI4DMAIl00l
;
reg
CAXI4DMAll00l
;
localparam
[
7
:
0
]
CAXI4DMAO1OII
=
8
'b
00000001
;
localparam
[
7
:
0
]
CAXI4DMAO000l
=
8
'b
00000010
;
localparam
[
7
:
0
]
CAXI4DMAI000l
=
8
'b
00000100
;
localparam
[
7
:
0
]
CAXI4DMAl000l
=
8
'b
00001000
;
localparam
[
7
:
0
]
CAXI4DMAO100l
=
8
'b
00010000
;
localparam
[
7
:
0
]
CAXI4DMAI100l
=
8
'b
00100000
;
localparam
[
7
:
0
]
CAXI4DMAl100l
=
8
'b
01000000
;
localparam
[
7
:
0
]
CAXI4DMAOO10l
=
8
'b
10000000
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAOIl0l
<=
1
'b
0
;
CAXI4DMAlIl0l
<=
32
'b
0
;
CAXI4DMAIll0l
<=
1
'b
0
;
CAXI4DMAOOOl
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAO0l0l
<=
32
'b
0
;
CAXI4DMAl0l0l
<=
2
'b
0
;
CAXI4DMAI1l0l
<=
3
'b
0
;
CAXI4DMAOO00l
<=
1
'b
0
;
CAXI4DMAlO00l
<=
1
'b
0
;
CAXI4DMAIOl0l
<=
1
'b
0
;
CAXI4DMAlI0ll
<=
1
'b
0
;
CAXI4DMAII00l
<=
1
'b
0
;
CAXI4DMAOl00l
<=
{
CAXI4DMAI1OI
{
1
'b
0
}
}
;
CAXI4DMAll00l
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAOOOIl
)
begin
if
(
CAXI4DMAIOOIl
==
2
'b
00
)
begin
CAXI4DMAOO00l
<=
1
'b
1
;
CAXI4DMAlO00l
<=
1
'b
1
;
CAXI4DMAll00l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO10l
;
end
else
if
(
CAXI4DMAII0OI
)
begin
if
(
CAXI4DMAI0OIl
)
begin
CAXI4DMAIll0l
<=
1
'b
1
;
CAXI4DMAO0l0l
<=
CAXI4DMAIIOIl
;
CAXI4DMAl0l0l
<=
CAXI4DMAIOOIl
;
CAXI4DMAI1l0l
<=
CAXI4DMAlOOIl
;
CAXI4DMAOOOl
<=
CAXI4DMAlIOIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAl100l
;
if
(
CAXI4DMAllllI
==
8
'b
00000001
)
begin
CAXI4DMAOl00l
<=
PRI_0_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000010
)
begin
CAXI4DMAOl00l
<=
PRI_1_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000100
)
begin
CAXI4DMAOl00l
<=
PRI_2_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00001000
)
begin
CAXI4DMAOl00l
<=
PRI_3_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00010000
)
begin
CAXI4DMAOl00l
<=
PRI_4_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00100000
)
begin
CAXI4DMAOl00l
<=
PRI_5_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
01000000
)
begin
CAXI4DMAOl00l
<=
PRI_6_NUM_OF_BEATS
;
end
else
begin
CAXI4DMAOl00l
<=
PRI_7_NUM_OF_BEATS
;
end
end
else
begin
CAXI4DMAOIl0l
<=
1
'b
1
;
CAXI4DMAlIl0l
<=
CAXI4DMAlI0OI
;
CAXI4DMAOO1OI
<=
CAXI4DMAO000l
;
end
end
else
begin
CAXI4DMAIll0l
<=
1
'b
1
;
CAXI4DMAO0l0l
<=
CAXI4DMAIIOIl
;
CAXI4DMAl0l0l
<=
CAXI4DMAIOOIl
;
CAXI4DMAI1l0l
<=
CAXI4DMAlOOIl
;
CAXI4DMAOOOl
<=
CAXI4DMAlIOIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAl100l
;
if
(
CAXI4DMAllllI
==
8
'b
00000001
)
begin
CAXI4DMAOl00l
<=
PRI_0_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000010
)
begin
CAXI4DMAOl00l
<=
PRI_1_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000100
)
begin
CAXI4DMAOl00l
<=
PRI_2_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00001000
)
begin
CAXI4DMAOl00l
<=
PRI_3_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00010000
)
begin
CAXI4DMAOl00l
<=
PRI_4_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00100000
)
begin
CAXI4DMAOl00l
<=
PRI_5_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
01000000
)
begin
CAXI4DMAOl00l
<=
PRI_6_NUM_OF_BEATS
;
end
else
begin
CAXI4DMAOl00l
<=
PRI_7_NUM_OF_BEATS
;
end
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAOO10l
:
begin
if
(
CAXI4DMAl10Ol
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAll00l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO10l
;
end
end
CAXI4DMAO000l
:
begin
if
(
CAXI4DMAlII1I
)
begin
if
(
CAXI4DMAOlI1I
)
begin
CAXI4DMAIll0l
<=
1
'b
1
;
CAXI4DMAO0l0l
<=
CAXI4DMAIIOIl
;
CAXI4DMAl0l0l
<=
CAXI4DMAIOOIl
;
CAXI4DMAI1l0l
<=
CAXI4DMAlOOIl
;
CAXI4DMAOOOl
<=
CAXI4DMAlIOIl
;
if
(
CAXI4DMAllllI
==
8
'b
00000001
)
begin
CAXI4DMAOl00l
<=
PRI_0_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000010
)
begin
CAXI4DMAOl00l
<=
PRI_1_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000100
)
begin
CAXI4DMAOl00l
<=
PRI_2_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00001000
)
begin
CAXI4DMAOl00l
<=
PRI_3_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00010000
)
begin
CAXI4DMAOl00l
<=
PRI_4_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00100000
)
begin
CAXI4DMAOl00l
<=
PRI_5_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
01000000
)
begin
CAXI4DMAOl00l
<=
PRI_6_NUM_OF_BEATS
;
end
else
begin
CAXI4DMAOl00l
<=
PRI_7_NUM_OF_BEATS
;
end
if
(
CAXI4DMAl011
)
begin
CAXI4DMAOO00l
<=
1
'b
1
;
CAXI4DMAlO00l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI000l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl100l
;
end
end
else
begin
CAXI4DMAOO00l
<=
1
'b
1
;
CAXI4DMAII00l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI100l
;
end
end
else
begin
CAXI4DMAOIl0l
<=
1
'b
1
;
CAXI4DMAlIl0l
<=
CAXI4DMAlI0OI
;
CAXI4DMAOO1OI
<=
CAXI4DMAO000l
;
end
end
CAXI4DMAl100l
:
begin
if
(
CAXI4DMAl011
)
begin
CAXI4DMAOO00l
<=
1
'b
1
;
CAXI4DMAlO00l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI000l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl100l
;
end
end
CAXI4DMAI000l
:
begin
if
(
CAXI4DMAl0OIl
)
begin
CAXI4DMAIOl0l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAl000l
;
end
else
if
(
CAXI4DMAO1OIl
)
begin
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO100l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAI000l
;
end
end
CAXI4DMAl000l
:
begin
if
(
CAXI4DMAI1OIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAIOl0l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAl000l
;
end
end
CAXI4DMAO100l
:
begin
if
(
CAXI4DMAl1OIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO100l
;
end
end
CAXI4DMAI100l
:
begin
if
(
CAXI4DMAOlIOl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAII00l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI100l
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOOl0l
<=
1
'b
0
;
end
else
begin
CAXI4DMAOOl0l
<=
CAXI4DMAIOl0l
;
end
end
assign
CAXI4DMAOOIIl
=
CAXI4DMAOOl0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAII0ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAII0ll
<=
CAXI4DMAlI0ll
;
end
end
assign
CAXI4DMAIllOI
=
CAXI4DMAII0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlOl0l
<=
1
'b
0
;
end
else
begin
CAXI4DMAlOl0l
<=
CAXI4DMAOIl0l
;
end
end
assign
CAXI4DMAO1O1I
=
CAXI4DMAlOl0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIIl0l
<=
32
'b
0
;
end
else
begin
CAXI4DMAIIl0l
<=
CAXI4DMAlIl0l
;
end
end
assign
CAXI4DMAOIl0I
=
CAXI4DMAIIl0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOll0l
<=
1
'b
0
;
end
else
begin
CAXI4DMAOll0l
<=
CAXI4DMAIll0l
;
end
end
assign
CAXI4DMAII
=
CAXI4DMAOll0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl11I
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAl11I
<=
CAXI4DMAOOOl
;
end
end
assign
CAXI4DMAOl
=
CAXI4DMAl11I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlll0l
<=
32
'b
0
;
end
else
begin
CAXI4DMAlll0l
<=
CAXI4DMAO0l0l
;
end
end
assign
CAXI4DMAO101I
=
CAXI4DMAlll0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI0l0l
<=
2
'b
0
;
end
else
begin
CAXI4DMAI0l0l
<=
CAXI4DMAl0l0l
;
end
end
assign
CAXI4DMAlI
=
CAXI4DMAI0l0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO1l0l
<=
3
'b
0
;
end
else
begin
CAXI4DMAO1l0l
<=
CAXI4DMAI1l0l
;
end
end
assign
CAXI4DMAll
=
CAXI4DMAO1l0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl1l0l
<=
1
'b
0
;
end
else
begin
CAXI4DMAl1l0l
<=
CAXI4DMAOO00l
;
end
end
assign
CAXI4DMAlOlOl
=
CAXI4DMAl1l0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO00l
<=
1
'b
0
;
end
else
begin
CAXI4DMAIO00l
<=
CAXI4DMAlO00l
;
end
end
assign
CAXI4DMAIIllI
=
CAXI4DMAIO00l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOI00l
<=
1
'b
0
;
end
else
begin
CAXI4DMAOI00l
<=
CAXI4DMAII00l
;
end
end
assign
CAXI4DMAO1OOl
=
CAXI4DMAOI00l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI00l
<=
{
CAXI4DMAI1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAlI00l
<=
CAXI4DMAOl00l
;
end
end
assign
CAXI4DMAO0
=
CAXI4DMAlI00l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIl00l
<=
1
'b
0
;
end
else
begin
CAXI4DMAIl00l
<=
CAXI4DMAll00l
;
end
end
assign
CAXI4DMAO10Ol
=
CAXI4DMAIl00l
;
endmodule
