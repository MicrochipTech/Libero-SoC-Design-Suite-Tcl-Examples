`timescale 1ns / 1ns
///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: MICROSEMI
//
// IP Core: COREAXI4INTERCONNECT
//
//  Description  : The AMBA AXI4 Interconnect core connects one or more AXI memory-mapped master devices to one or
//                 more memory-mapped slave devices. The AMBA AXI protocol supports high-performance, high-frequency
//                 system designs. This file provides an AXI4Interconnect between up to 8 masters and 32 slaves. 
//                 All ports Master buses can be AHB-Lite, AXI3, AXI4 or AXI4-Lite and all ports Slave buses can be 
//                 AXI3, AXI4 or AXI4-Lite Infrastructure components ensure all ports are converted to AXI4 to be 
//                 switched by caxi4interconnect_Axi4CrossBar.
//                                                               
//                 Note: AXI3 Interleaving not supported in AXI3 interface module. 
//
//  COPYRIGHT 2017 BY MICROSEMI 
//  THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
//  FROM MICROSEMI CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
//  MICROSEMI FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
//  NO BACK-UP OF THE FILE SHOULD BE MADE. 
//
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

module COREAXI4INTERCONNECT

  (
  
   // Global Signals
  ACLK,
  ARESETN,

  M_CLK0,
  M_CLK1,
  M_CLK2,
  M_CLK3,
  M_CLK4,
  M_CLK5,
  M_CLK6,
  M_CLK7,

  S_CLK0,
  S_CLK1,
  S_CLK2,
  S_CLK3,
  S_CLK4,
  S_CLK5,
  S_CLK6,
  S_CLK7,

// Expansion to 32 slave ports  
  S_CLK8,
  S_CLK9,
  S_CLK10,
  S_CLK11,
  S_CLK12,
  S_CLK13,
  S_CLK14,
  S_CLK15,
  S_CLK16,
  S_CLK17,
  S_CLK18,
  S_CLK19,
  S_CLK20,
  S_CLK21,
  S_CLK22,
  S_CLK23,
  S_CLK24,
  S_CLK25,
  S_CLK26,
  S_CLK27,
  S_CLK28,
  S_CLK29,
  S_CLK30,
  S_CLK31,

   // Master Write Address Ports
  MASTER0_AWID,
  MASTER0_AWADDR,
  MASTER0_AWLEN,
  MASTER0_AWSIZE,
  MASTER0_AWBURST,
  MASTER0_AWLOCK,
  MASTER0_AWCACHE,
  MASTER0_AWPROT,
  MASTER0_AWREGION,
  MASTER0_AWQOS,        // not used internally
  MASTER0_AWUSER,        // not used internally
  MASTER0_AWVALID,
  MASTER0_AWREADY,

  MASTER1_AWID,
  MASTER1_AWADDR,
  MASTER1_AWLEN,
  MASTER1_AWSIZE,
  MASTER1_AWBURST,
  MASTER1_AWLOCK,
  MASTER1_AWCACHE,
  MASTER1_AWPROT,
  MASTER1_AWREGION,
  MASTER1_AWQOS,        // not used internally
  MASTER1_AWUSER,        // not used internally
  MASTER1_AWVALID,
  MASTER1_AWREADY,

  MASTER2_AWID,
  MASTER2_AWADDR,
  MASTER2_AWLEN,
  MASTER2_AWSIZE,
  MASTER2_AWBURST,
  MASTER2_AWLOCK,
  MASTER2_AWCACHE,
  MASTER2_AWPROT,
  MASTER2_AWREGION,
  MASTER2_AWQOS,        // not used internally
  MASTER2_AWUSER,        // not used internally
  MASTER2_AWVALID,
  MASTER2_AWREADY,  

  MASTER3_AWID,
  MASTER3_AWADDR,
  MASTER3_AWLEN,
  MASTER3_AWSIZE,
  MASTER3_AWBURST,
  MASTER3_AWLOCK,
  MASTER3_AWCACHE,
  MASTER3_AWPROT,
  MASTER3_AWREGION,
  MASTER3_AWQOS,        // not used internally
  MASTER3_AWUSER,        // not used internally
  MASTER3_AWVALID,
  MASTER3_AWREADY,    
  
  MASTER4_AWID,
  MASTER4_AWADDR,
  MASTER4_AWLEN,
  MASTER4_AWSIZE,
  MASTER4_AWBURST,
  MASTER4_AWLOCK,
  MASTER4_AWCACHE,
  MASTER4_AWPROT,
  MASTER4_AWREGION,
  MASTER4_AWQOS,        // not used internally
  MASTER4_AWUSER,        // not used internally
  MASTER4_AWVALID,
  MASTER4_AWREADY,    
  
  MASTER5_AWID,
  MASTER5_AWADDR,
  MASTER5_AWLEN,
  MASTER5_AWSIZE,
  MASTER5_AWBURST,
  MASTER5_AWLOCK,
  MASTER5_AWCACHE,
  MASTER5_AWPROT,
  MASTER5_AWREGION,
  MASTER5_AWQOS,        // not used internally
  MASTER5_AWUSER,        // not used internally
  MASTER5_AWVALID,
  MASTER5_AWREADY,
  
  MASTER6_AWID,
  MASTER6_AWADDR,
  MASTER6_AWLEN,
  MASTER6_AWSIZE,
  MASTER6_AWBURST,
  MASTER6_AWLOCK,
  MASTER6_AWCACHE,
  MASTER6_AWPROT,
  MASTER6_AWREGION,
  MASTER6_AWQOS,        // not used internally
  MASTER6_AWUSER,        // not used internally
  MASTER6_AWVALID,
  MASTER6_AWREADY,  

  MASTER7_AWID,
  MASTER7_AWADDR,
  MASTER7_AWLEN,
  MASTER7_AWSIZE,
  MASTER7_AWBURST,
  MASTER7_AWLOCK,
  MASTER7_AWCACHE,
  MASTER7_AWPROT,
  MASTER7_AWREGION,
  MASTER7_AWQOS,        // not used internally
  MASTER7_AWUSER,        // not used internally
  MASTER7_AWVALID,
  MASTER7_AWREADY,  
  
   // Master Write Data Ports
  MASTER0_WDATA,
  MASTER0_WSTRB,
  MASTER0_WLAST,
  MASTER0_WUSER,
  MASTER0_WVALID,
  MASTER0_WREADY,
 
   MASTER1_WDATA,
  MASTER1_WSTRB,
  MASTER1_WLAST,
  MASTER1_WUSER,
  MASTER1_WVALID,
  MASTER1_WREADY,
 
   MASTER2_WDATA,
  MASTER2_WSTRB,
  MASTER2_WLAST,
  MASTER2_WUSER,
  MASTER2_WVALID,
  MASTER2_WREADY,
 
   MASTER3_WDATA,
  MASTER3_WSTRB,
  MASTER3_WLAST,
  MASTER3_WUSER,
  MASTER3_WVALID,
  MASTER3_WREADY,
  
  MASTER4_WDATA,
  MASTER4_WSTRB,
  MASTER4_WLAST,
  MASTER4_WUSER,
  MASTER4_WVALID,
  MASTER4_WREADY,
  
  MASTER5_WDATA,
  MASTER5_WSTRB,
  MASTER5_WLAST,
  MASTER5_WUSER,
  MASTER5_WVALID,
  MASTER5_WREADY,
  
  MASTER6_WDATA,
  MASTER6_WSTRB,
  MASTER6_WLAST,
  MASTER6_WUSER,
  MASTER6_WVALID,
  MASTER6_WREADY,
  
  MASTER7_WDATA,
  MASTER7_WSTRB,
  MASTER7_WLAST,
  MASTER7_WUSER,
  MASTER7_WVALID,
  MASTER7_WREADY,
  
  // Master Write Response Ports
  MASTER0_BID,
  MASTER0_BRESP,
  MASTER0_BUSER,
  MASTER0_BVALID,
  MASTER0_BREADY,

  MASTER1_BID,
  MASTER1_BRESP,
  MASTER1_BUSER,
  MASTER1_BVALID,
  MASTER1_BREADY,  
  
  MASTER2_BID,
  MASTER2_BRESP,
  MASTER2_BUSER,
  MASTER2_BVALID,
  MASTER2_BREADY,  

  MASTER3_BID,
  MASTER3_BRESP,
  MASTER3_BUSER,
  MASTER3_BVALID,
  MASTER3_BREADY,  
  
  MASTER4_BID,
  MASTER4_BRESP,
  MASTER4_BUSER,
  MASTER4_BVALID,
  MASTER4_BREADY,  
  
  MASTER5_BID,
  MASTER5_BRESP,
  MASTER5_BUSER,
  MASTER5_BVALID,
  MASTER5_BREADY,  
  
  MASTER6_BID,
  MASTER6_BRESP,
  MASTER6_BUSER,
  MASTER6_BVALID,
  MASTER6_BREADY,  
  
  MASTER7_BID,
  MASTER7_BRESP,
  MASTER7_BUSER,
  MASTER7_BVALID,
  MASTER7_BREADY,  
  
   // Master Read Address Ports
  MASTER0_ARID,
  MASTER0_ARADDR,
  MASTER0_ARLEN,
  MASTER0_ARSIZE,
  MASTER0_ARBURST,
  MASTER0_ARLOCK,
  MASTER0_ARCACHE,
  MASTER0_ARPROT,
  MASTER0_ARREGION,
  MASTER0_ARQOS,    // not used
  MASTER0_ARUSER,
  MASTER0_ARVALID,
  MASTER0_ARREADY,
  
  MASTER1_ARID,
  MASTER1_ARADDR,
  MASTER1_ARLEN,
  MASTER1_ARSIZE,
  MASTER1_ARBURST,
  MASTER1_ARLOCK,
  MASTER1_ARCACHE,
  MASTER1_ARPROT,
  MASTER1_ARREGION,
  MASTER1_ARQOS,    // not used
  MASTER1_ARUSER,
  MASTER1_ARVALID,
  MASTER1_ARREADY,  

  MASTER2_ARID,
  MASTER2_ARADDR,
  MASTER2_ARLEN,
  MASTER2_ARSIZE,
  MASTER2_ARBURST,
  MASTER2_ARLOCK,
  MASTER2_ARCACHE,
  MASTER2_ARPROT,
  MASTER2_ARREGION,
  MASTER2_ARQOS,    // not used
  MASTER2_ARUSER,
  MASTER2_ARVALID,
  MASTER2_ARREADY,  
  
  MASTER3_ARID,
  MASTER3_ARADDR,
  MASTER3_ARLEN,
  MASTER3_ARSIZE,
  MASTER3_ARBURST,
  MASTER3_ARLOCK,
  MASTER3_ARCACHE,
  MASTER3_ARPROT,
  MASTER3_ARREGION,
  MASTER3_ARQOS,    // not used
  MASTER3_ARUSER,
  MASTER3_ARVALID,
  MASTER3_ARREADY,  
  
  MASTER4_ARID,
  MASTER4_ARADDR,
  MASTER4_ARLEN,
  MASTER4_ARSIZE,
  MASTER4_ARBURST,
  MASTER4_ARLOCK,
  MASTER4_ARCACHE,
  MASTER4_ARPROT,
  MASTER4_ARREGION,
  MASTER4_ARQOS,    // not used
  MASTER4_ARUSER,
  MASTER4_ARVALID,
  MASTER4_ARREADY,  
  
  MASTER5_ARID,
  MASTER5_ARADDR,
  MASTER5_ARLEN,
  MASTER5_ARSIZE,
  MASTER5_ARBURST,
  MASTER5_ARLOCK,
  MASTER5_ARCACHE,
  MASTER5_ARPROT,
  MASTER5_ARREGION,
  MASTER5_ARQOS,    // not used
  MASTER5_ARUSER,
  MASTER5_ARVALID,
  MASTER5_ARREADY,  
  
  MASTER6_ARID,
  MASTER6_ARADDR,
  MASTER6_ARLEN,
  MASTER6_ARSIZE,
  MASTER6_ARBURST,
  MASTER6_ARLOCK,
  MASTER6_ARCACHE,
  MASTER6_ARPROT,
  MASTER6_ARREGION,
  MASTER6_ARQOS,    // not used
  MASTER6_ARUSER,
  MASTER6_ARVALID,
  MASTER6_ARREADY,  
  
  MASTER7_ARID,
  MASTER7_ARADDR,
  MASTER7_ARLEN,
  MASTER7_ARSIZE,
  MASTER7_ARBURST,
  MASTER7_ARLOCK,
  MASTER7_ARCACHE,
  MASTER7_ARPROT,
  MASTER7_ARREGION,
  MASTER7_ARQOS,    // not used
  MASTER7_ARUSER,
  MASTER7_ARVALID,
  MASTER7_ARREADY,  
  
   // Master Read Data Ports
  MASTER0_RID,
  MASTER0_RDATA,
  MASTER0_RRESP,
  MASTER0_RLAST,
  MASTER0_RUSER,
  MASTER0_RVALID,
  MASTER0_RREADY,
 
  MASTER1_RID,
  MASTER1_RDATA,
  MASTER1_RRESP,
  MASTER1_RLAST,
  MASTER1_RUSER,
  MASTER1_RVALID,
  MASTER1_RREADY,
   
  MASTER2_RID,
  MASTER2_RDATA,
  MASTER2_RRESP,
  MASTER2_RLAST,
  MASTER2_RUSER,
  MASTER2_RVALID,
  MASTER2_RREADY,
   
  MASTER3_RID,
  MASTER3_RDATA,
  MASTER3_RRESP,
  MASTER3_RLAST,
  MASTER3_RUSER,
  MASTER3_RVALID,
  MASTER3_RREADY,
  
  MASTER4_RID,
  MASTER4_RDATA,
  MASTER4_RRESP,
  MASTER4_RLAST,
  MASTER4_RUSER,
  MASTER4_RVALID,
  MASTER4_RREADY,
  
  MASTER5_RID,
  MASTER5_RDATA,
  MASTER5_RRESP,
  MASTER5_RLAST,
  MASTER5_RUSER,
  MASTER5_RVALID,
  MASTER5_RREADY,
  
  MASTER6_RID,
  MASTER6_RDATA,
  MASTER6_RRESP,
  MASTER6_RLAST,
  MASTER6_RUSER,
  MASTER6_RVALID,
  MASTER6_RREADY,
  
  MASTER7_RID,
  MASTER7_RDATA,
  MASTER7_RRESP,
  MASTER7_RLAST,
  MASTER7_RUSER,
  MASTER7_RVALID,
  MASTER7_RREADY,
      
  // AHB Masters
   MASTER0_HADDR,
  MASTER0_HBURST,
  MASTER0_HMASTLOCK,
  MASTER0_HPROT,          
  MASTER0_HSIZE,
  MASTER0_HNONSEC,
  MASTER0_HTRANS,
  MASTER0_HWDATA,
  MASTER0_HRDATA,
  MASTER0_HWRITE,
  MASTER0_HREADY,
  MASTER0_HRESP,
//  MASTER0_HEXOKAY,
//  MASTER0_HEXCL,
  MASTER0_HSEL,

  MASTER1_HADDR,
  MASTER1_HBURST,
  MASTER1_HMASTLOCK,
  MASTER1_HPROT,          
  MASTER1_HSIZE,
  MASTER1_HNONSEC,
  MASTER1_HTRANS,
  MASTER1_HWDATA,
  MASTER1_HRDATA,
  MASTER1_HWRITE,
  MASTER1_HREADY,
  MASTER1_HRESP,
//  MASTER1_HEXOKAY,
//  MASTER1_HEXCL,
  MASTER1_HSEL,

  MASTER2_HADDR,
  MASTER2_HBURST,
  MASTER2_HMASTLOCK,
  MASTER2_HPROT,          
  MASTER2_HSIZE,
  MASTER2_HNONSEC,
  MASTER2_HTRANS,
  MASTER2_HWDATA,
  MASTER2_HRDATA,
  MASTER2_HWRITE,
  MASTER2_HREADY,
  MASTER2_HRESP,
//  MASTER2_HEXOKAY,
//  MASTER2_HEXCL,
  MASTER2_HSEL,

  MASTER3_HADDR,
  MASTER3_HBURST,
  MASTER3_HMASTLOCK,
  MASTER3_HPROT,          
  MASTER3_HSIZE,
  MASTER3_HNONSEC,
  MASTER3_HTRANS,
  MASTER3_HWDATA,
  MASTER3_HRDATA,
  MASTER3_HWRITE,
  MASTER3_HREADY,
  MASTER3_HRESP,
//  MASTER3_HEXOKAY,
//  MASTER3_HEXCL,
  MASTER3_HSEL,

  MASTER4_HADDR,
  MASTER4_HBURST,
  MASTER4_HMASTLOCK,
  MASTER4_HPROT,          
  MASTER4_HSIZE,
  MASTER4_HNONSEC,
  MASTER4_HTRANS,
  MASTER4_HWDATA,
  MASTER4_HRDATA,
  MASTER4_HWRITE,
  MASTER4_HREADY,
  MASTER4_HRESP,
//  MASTER4_HEXOKAY,
//  MASTER4_HEXCL,
  MASTER4_HSEL,

  MASTER5_HADDR,
  MASTER5_HBURST,
  MASTER5_HMASTLOCK,
  MASTER5_HPROT,          
  MASTER5_HSIZE,
  MASTER5_HNONSEC,
  MASTER5_HTRANS,
  MASTER5_HWDATA,
  MASTER5_HRDATA,
  MASTER5_HWRITE,
  MASTER5_HREADY,
  MASTER5_HRESP,
//  MASTER5_HEXOKAY,
//  MASTER5_HEXCL,
  MASTER5_HSEL,

  MASTER6_HADDR,
  MASTER6_HBURST,
  MASTER6_HMASTLOCK,
  MASTER6_HPROT,          
  MASTER6_HSIZE,
  MASTER6_HNONSEC,
  MASTER6_HTRANS,
  MASTER6_HWDATA,
  MASTER6_HRDATA,
  MASTER6_HWRITE,
  MASTER6_HREADY,
  MASTER6_HRESP,
//  MASTER6_HEXOKAY,
//  MASTER6_HEXCL,
  MASTER6_HSEL,

  MASTER7_HADDR,
  MASTER7_HBURST,
  MASTER7_HMASTLOCK,
  MASTER7_HPROT,          
  MASTER7_HSIZE,
  MASTER7_HNONSEC,
  MASTER7_HTRANS,
  MASTER7_HWDATA,
  MASTER7_HRDATA,
  MASTER7_HWRITE,
  MASTER7_HREADY,
  MASTER7_HRESP,
//  MASTER7_HEXOKAY,
//  MASTER7_HEXCL,
  MASTER7_HSEL,

  // Slave Write Address Port
  SLAVE0_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE0_AWADDR,
  SLAVE0_AWLEN,
  SLAVE0_AWSIZE,
  SLAVE0_AWBURST,
  SLAVE0_AWLOCK,
  SLAVE0_AWCACHE,
  SLAVE0_AWPROT,
  SLAVE0_AWREGION,    // not used
  SLAVE0_AWQOS,      // not used
  SLAVE0_AWUSER,
  SLAVE0_AWVALID,
  SLAVE0_AWREADY,
  
  SLAVE1_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE1_AWADDR,
  SLAVE1_AWLEN,
  SLAVE1_AWSIZE,
  SLAVE1_AWBURST,
  SLAVE1_AWLOCK,
  SLAVE1_AWCACHE,
  SLAVE1_AWPROT,
  SLAVE1_AWREGION,    // not used
  SLAVE1_AWQOS,      // not used
  SLAVE1_AWUSER,
  SLAVE1_AWVALID,
  SLAVE1_AWREADY,  
 
  SLAVE2_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE2_AWADDR,
  SLAVE2_AWLEN,
  SLAVE2_AWSIZE,
  SLAVE2_AWBURST,
  SLAVE2_AWLOCK,
  SLAVE2_AWCACHE,
  SLAVE2_AWPROT,
  SLAVE2_AWREGION,    // not used
  SLAVE2_AWQOS,      // not used
  SLAVE2_AWUSER,
  SLAVE2_AWVALID,
  SLAVE2_AWREADY, 
   
  SLAVE3_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE3_AWADDR,
  SLAVE3_AWLEN,
  SLAVE3_AWSIZE,
  SLAVE3_AWBURST,
  SLAVE3_AWLOCK,
  SLAVE3_AWCACHE,
  SLAVE3_AWPROT,
  SLAVE3_AWREGION,    // not used
  SLAVE3_AWQOS,      // not used
  SLAVE3_AWUSER,
  SLAVE3_AWVALID,
  SLAVE3_AWREADY,

  SLAVE4_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE4_AWADDR,
  SLAVE4_AWLEN,
  SLAVE4_AWSIZE,
  SLAVE4_AWBURST,
  SLAVE4_AWLOCK,
  SLAVE4_AWCACHE,
  SLAVE4_AWPROT,
  SLAVE4_AWREGION,    // not used
  SLAVE4_AWQOS,      // not used
  SLAVE4_AWUSER,
  SLAVE4_AWVALID,
  SLAVE4_AWREADY,
  
  SLAVE5_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE5_AWADDR,
  SLAVE5_AWLEN,
  SLAVE5_AWSIZE,
  SLAVE5_AWBURST,
  SLAVE5_AWLOCK,
  SLAVE5_AWCACHE,
  SLAVE5_AWPROT,
  SLAVE5_AWREGION,    // not used
  SLAVE5_AWQOS,      // not used
  SLAVE5_AWUSER,
  SLAVE5_AWVALID,
  SLAVE5_AWREADY,  

  SLAVE6_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE6_AWADDR,
  SLAVE6_AWLEN,
  SLAVE6_AWSIZE,
  SLAVE6_AWBURST,
  SLAVE6_AWLOCK,
  SLAVE6_AWCACHE,
  SLAVE6_AWPROT,
  SLAVE6_AWREGION,    // not used
  SLAVE6_AWQOS,      // not used
  SLAVE6_AWUSER,
  SLAVE6_AWVALID,
  SLAVE6_AWREADY,  
  
  SLAVE7_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE7_AWADDR,
  SLAVE7_AWLEN,
  SLAVE7_AWSIZE,
  SLAVE7_AWBURST,
  SLAVE7_AWLOCK,
  SLAVE7_AWCACHE,
  SLAVE7_AWPROT,
  SLAVE7_AWREGION,    // not used
  SLAVE7_AWQOS,      // not used
  SLAVE7_AWUSER,
  SLAVE7_AWVALID,
  SLAVE7_AWREADY,
  
  SLAVE8_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE8_AWADDR,
  SLAVE8_AWLEN,
  SLAVE8_AWSIZE,
  SLAVE8_AWBURST,
  SLAVE8_AWLOCK,
  SLAVE8_AWCACHE,
  SLAVE8_AWPROT,
  SLAVE8_AWREGION,    // not used
  SLAVE8_AWQOS,      // not used
  SLAVE8_AWUSER,
  SLAVE8_AWVALID,
  SLAVE8_AWREADY,  
  
  SLAVE9_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE9_AWADDR,
  SLAVE9_AWLEN,
  SLAVE9_AWSIZE,
  SLAVE9_AWBURST,
  SLAVE9_AWLOCK,
  SLAVE9_AWCACHE,
  SLAVE9_AWPROT,
  SLAVE9_AWREGION,    // not used
  SLAVE9_AWQOS,      // not used
  SLAVE9_AWUSER,
  SLAVE9_AWVALID,
  SLAVE9_AWREADY,  
  
  SLAVE10_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE10_AWADDR,
  SLAVE10_AWLEN,
  SLAVE10_AWSIZE,
  SLAVE10_AWBURST,
  SLAVE10_AWLOCK,
  SLAVE10_AWCACHE,
  SLAVE10_AWPROT,
  SLAVE10_AWREGION,    // not used
  SLAVE10_AWQOS,      // not used
  SLAVE10_AWUSER,
  SLAVE10_AWVALID,
  SLAVE10_AWREADY,  
  
  SLAVE11_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE11_AWADDR,
  SLAVE11_AWLEN,
  SLAVE11_AWSIZE,
  SLAVE11_AWBURST,
  SLAVE11_AWLOCK,
  SLAVE11_AWCACHE,
  SLAVE11_AWPROT,
  SLAVE11_AWREGION,    // not used
  SLAVE11_AWQOS,      // not used
  SLAVE11_AWUSER,
  SLAVE11_AWVALID,
  SLAVE11_AWREADY,  
   
  SLAVE12_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE12_AWADDR,
  SLAVE12_AWLEN,
  SLAVE12_AWSIZE,
  SLAVE12_AWBURST,
  SLAVE12_AWLOCK,
  SLAVE12_AWCACHE,
  SLAVE12_AWPROT,
  SLAVE12_AWREGION,    // not used
  SLAVE12_AWQOS,      // not used
  SLAVE12_AWUSER,
  SLAVE12_AWVALID,
  SLAVE12_AWREADY,  
  
  SLAVE13_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE13_AWADDR,
  SLAVE13_AWLEN,
  SLAVE13_AWSIZE,
  SLAVE13_AWBURST,
  SLAVE13_AWLOCK,
  SLAVE13_AWCACHE,
  SLAVE13_AWPROT,
  SLAVE13_AWREGION,    // not used
  SLAVE13_AWQOS,      // not used
  SLAVE13_AWUSER,
  SLAVE13_AWVALID,
  SLAVE13_AWREADY,  
  
  SLAVE14_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE14_AWADDR,
  SLAVE14_AWLEN,
  SLAVE14_AWSIZE,
  SLAVE14_AWBURST,
  SLAVE14_AWLOCK,
  SLAVE14_AWCACHE,
  SLAVE14_AWPROT,
  SLAVE14_AWREGION,    // not used
  SLAVE14_AWQOS,      // not used
  SLAVE14_AWUSER,
  SLAVE14_AWVALID,
  SLAVE14_AWREADY,  
  
  SLAVE15_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE15_AWADDR,
  SLAVE15_AWLEN,
  SLAVE15_AWSIZE,
  SLAVE15_AWBURST,
  SLAVE15_AWLOCK,
  SLAVE15_AWCACHE,
  SLAVE15_AWPROT,
  SLAVE15_AWREGION,    // not used
  SLAVE15_AWQOS,      // not used
  SLAVE15_AWUSER,
  SLAVE15_AWVALID,
  SLAVE15_AWREADY,  
  
  SLAVE16_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE16_AWADDR,
  SLAVE16_AWLEN,
  SLAVE16_AWSIZE,
  SLAVE16_AWBURST,
  SLAVE16_AWLOCK,
  SLAVE16_AWCACHE,
  SLAVE16_AWPROT,
  SLAVE16_AWREGION,    // not used
  SLAVE16_AWQOS,      // not used
  SLAVE16_AWUSER,
  SLAVE16_AWVALID,
  SLAVE16_AWREADY,  
  
  SLAVE17_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE17_AWADDR,
  SLAVE17_AWLEN,
  SLAVE17_AWSIZE,
  SLAVE17_AWBURST,
  SLAVE17_AWLOCK,
  SLAVE17_AWCACHE,
  SLAVE17_AWPROT,
  SLAVE17_AWREGION,    // not used
  SLAVE17_AWQOS,      // not used
  SLAVE17_AWUSER,
  SLAVE17_AWVALID,
  SLAVE17_AWREADY,  
  
  SLAVE18_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE18_AWADDR,
  SLAVE18_AWLEN,
  SLAVE18_AWSIZE,
  SLAVE18_AWBURST,
  SLAVE18_AWLOCK,
  SLAVE18_AWCACHE,
  SLAVE18_AWPROT,
  SLAVE18_AWREGION,    // not used
  SLAVE18_AWQOS,      // not used
  SLAVE18_AWUSER,
  SLAVE18_AWVALID,
  SLAVE18_AWREADY,  
  
  SLAVE19_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE19_AWADDR,
  SLAVE19_AWLEN,
  SLAVE19_AWSIZE,
  SLAVE19_AWBURST,
  SLAVE19_AWLOCK,
  SLAVE19_AWCACHE,
  SLAVE19_AWPROT,
  SLAVE19_AWREGION,    // not used
  SLAVE19_AWQOS,      // not used
  SLAVE19_AWUSER,
  SLAVE19_AWVALID,
  SLAVE19_AWREADY,  
  
  SLAVE20_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE20_AWADDR,
  SLAVE20_AWLEN,
  SLAVE20_AWSIZE,
  SLAVE20_AWBURST,
  SLAVE20_AWLOCK,
  SLAVE20_AWCACHE,
  SLAVE20_AWPROT,
  SLAVE20_AWREGION,    // not used
  SLAVE20_AWQOS,      // not used
  SLAVE20_AWUSER,
  SLAVE20_AWVALID,
  SLAVE20_AWREADY,  
  
  SLAVE21_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE21_AWADDR,
  SLAVE21_AWLEN,
  SLAVE21_AWSIZE,
  SLAVE21_AWBURST,
  SLAVE21_AWLOCK,
  SLAVE21_AWCACHE,
  SLAVE21_AWPROT,
  SLAVE21_AWREGION,    // not used
  SLAVE21_AWQOS,      // not used
  SLAVE21_AWUSER,
  SLAVE21_AWVALID,
  SLAVE21_AWREADY,  
  
  SLAVE22_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE22_AWADDR,
  SLAVE22_AWLEN,
  SLAVE22_AWSIZE,
  SLAVE22_AWBURST,
  SLAVE22_AWLOCK,
  SLAVE22_AWCACHE,
  SLAVE22_AWPROT,
  SLAVE22_AWREGION,    // not used
  SLAVE22_AWQOS,      // not used
  SLAVE22_AWUSER,
  SLAVE22_AWVALID,
  SLAVE22_AWREADY,  
  
  SLAVE23_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE23_AWADDR,
  SLAVE23_AWLEN,
  SLAVE23_AWSIZE,
  SLAVE23_AWBURST,
  SLAVE23_AWLOCK,
  SLAVE23_AWCACHE,
  SLAVE23_AWPROT,
  SLAVE23_AWREGION,    // not used
  SLAVE23_AWQOS,      // not used
  SLAVE23_AWUSER,
  SLAVE23_AWVALID,
  SLAVE23_AWREADY,  
  
  SLAVE24_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE24_AWADDR,
  SLAVE24_AWLEN,
  SLAVE24_AWSIZE,
  SLAVE24_AWBURST,
  SLAVE24_AWLOCK,
  SLAVE24_AWCACHE,
  SLAVE24_AWPROT,
  SLAVE24_AWREGION,    // not used
  SLAVE24_AWQOS,      // not used
  SLAVE24_AWUSER,
  SLAVE24_AWVALID,
  SLAVE24_AWREADY,  
  
  SLAVE25_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE25_AWADDR,
  SLAVE25_AWLEN,
  SLAVE25_AWSIZE,
  SLAVE25_AWBURST,
  SLAVE25_AWLOCK,
  SLAVE25_AWCACHE,
  SLAVE25_AWPROT,
  SLAVE25_AWREGION,    // not used
  SLAVE25_AWQOS,      // not used
  SLAVE25_AWUSER,
  SLAVE25_AWVALID,
  SLAVE25_AWREADY,  
  
  SLAVE26_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE26_AWADDR,
  SLAVE26_AWLEN,
  SLAVE26_AWSIZE,
  SLAVE26_AWBURST,
  SLAVE26_AWLOCK,
  SLAVE26_AWCACHE,
  SLAVE26_AWPROT,
  SLAVE26_AWREGION,    // not used
  SLAVE26_AWQOS,      // not used
  SLAVE26_AWUSER,
  SLAVE26_AWVALID,
  SLAVE26_AWREADY,  
  
  SLAVE27_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE27_AWADDR,
  SLAVE27_AWLEN,
  SLAVE27_AWSIZE,
  SLAVE27_AWBURST,
  SLAVE27_AWLOCK,
  SLAVE27_AWCACHE,
  SLAVE27_AWPROT,
  SLAVE27_AWREGION,    // not used
  SLAVE27_AWQOS,      // not used
  SLAVE27_AWUSER,
  SLAVE27_AWVALID,
  SLAVE27_AWREADY,  
  
  SLAVE28_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE28_AWADDR,
  SLAVE28_AWLEN,
  SLAVE28_AWSIZE,
  SLAVE28_AWBURST,
  SLAVE28_AWLOCK,
  SLAVE28_AWCACHE,
  SLAVE28_AWPROT,
  SLAVE28_AWREGION,    // not used
  SLAVE28_AWQOS,      // not used
  SLAVE28_AWUSER,
  SLAVE28_AWVALID,
  SLAVE28_AWREADY,  
  
  SLAVE29_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE29_AWADDR,
  SLAVE29_AWLEN,
  SLAVE29_AWSIZE,
  SLAVE29_AWBURST,
  SLAVE29_AWLOCK,
  SLAVE29_AWCACHE,
  SLAVE29_AWPROT,
  SLAVE29_AWREGION,    // not used
  SLAVE29_AWQOS,      // not used
  SLAVE29_AWUSER,
  SLAVE29_AWVALID,
  SLAVE29_AWREADY,  
  
  SLAVE30_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE30_AWADDR,
  SLAVE30_AWLEN,
  SLAVE30_AWSIZE,
  SLAVE30_AWBURST,
  SLAVE30_AWLOCK,
  SLAVE30_AWCACHE,
  SLAVE30_AWPROT,
  SLAVE30_AWREGION,    // not used
  SLAVE30_AWQOS,      // not used
  SLAVE30_AWUSER,
  SLAVE30_AWVALID,
  SLAVE30_AWREADY,  
  
  SLAVE31_AWID,        // Slave ID is composed of Master Port ID concatenated with transaction ID
  SLAVE31_AWADDR,
  SLAVE31_AWLEN,
  SLAVE31_AWSIZE,
  SLAVE31_AWBURST,
  SLAVE31_AWLOCK,
  SLAVE31_AWCACHE,
  SLAVE31_AWPROT,
  SLAVE31_AWREGION,    // not used
  SLAVE31_AWQOS,      // not used
  SLAVE31_AWUSER,
  SLAVE31_AWVALID,
  SLAVE31_AWREADY,  
  
  
   // Slave Write Data Ports
  SLAVE0_WID,
  SLAVE0_WDATA,
  SLAVE0_WSTRB,
  SLAVE0_WLAST,
  SLAVE0_WUSER,
  SLAVE0_WVALID,
  SLAVE0_WREADY,

  SLAVE1_WID,
  SLAVE1_WDATA,
  SLAVE1_WSTRB,
  SLAVE1_WLAST,
  SLAVE1_WUSER,
  SLAVE1_WVALID,
  SLAVE1_WREADY,

  SLAVE2_WID,
  SLAVE2_WDATA,
  SLAVE2_WSTRB,
  SLAVE2_WLAST,
  SLAVE2_WUSER,
  SLAVE2_WVALID,
  SLAVE2_WREADY,  
  
  SLAVE3_WID,
  SLAVE3_WDATA,
  SLAVE3_WSTRB,
  SLAVE3_WLAST,
  SLAVE3_WUSER,
  SLAVE3_WVALID,
  SLAVE3_WREADY,  
  
  SLAVE4_WID,
  SLAVE4_WDATA,
  SLAVE4_WSTRB,
  SLAVE4_WLAST,
  SLAVE4_WUSER,
  SLAVE4_WVALID,
  SLAVE4_WREADY,  

  SLAVE5_WID,
  SLAVE5_WDATA,
  SLAVE5_WSTRB,
  SLAVE5_WLAST,
  SLAVE5_WUSER,
  SLAVE5_WVALID,
  SLAVE5_WREADY,  

  SLAVE6_WID,
  SLAVE6_WDATA,
  SLAVE6_WSTRB,
  SLAVE6_WLAST,
  SLAVE6_WUSER,
  SLAVE6_WVALID,
  SLAVE6_WREADY,

  SLAVE7_WID,
  SLAVE7_WDATA,
  SLAVE7_WSTRB,
  SLAVE7_WLAST,
  SLAVE7_WUSER,
  SLAVE7_WVALID,
  SLAVE7_WREADY,  

  SLAVE8_WID,
  SLAVE8_WDATA,
  SLAVE8_WSTRB,
  SLAVE8_WLAST,
  SLAVE8_WUSER,
  SLAVE8_WVALID,
  SLAVE8_WREADY,  

  SLAVE9_WID,
  SLAVE9_WDATA,
  SLAVE9_WSTRB,
  SLAVE9_WLAST,
  SLAVE9_WUSER,
  SLAVE9_WVALID,
  SLAVE9_WREADY,  

  SLAVE10_WID,
  SLAVE10_WDATA,
  SLAVE10_WSTRB,
  SLAVE10_WLAST,
  SLAVE10_WUSER,
  SLAVE10_WVALID,
  SLAVE10_WREADY,  

  SLAVE11_WID,
  SLAVE11_WDATA,
  SLAVE11_WSTRB,
  SLAVE11_WLAST,
  SLAVE11_WUSER,
  SLAVE11_WVALID,
  SLAVE11_WREADY,  

  SLAVE12_WID,
  SLAVE12_WDATA,
  SLAVE12_WSTRB,
  SLAVE12_WLAST,
  SLAVE12_WUSER,
  SLAVE12_WVALID,
  SLAVE12_WREADY,  

  SLAVE13_WID,
  SLAVE13_WDATA,
  SLAVE13_WSTRB,
  SLAVE13_WLAST,
  SLAVE13_WUSER,
  SLAVE13_WVALID,
  SLAVE13_WREADY,  

  SLAVE14_WID,
  SLAVE14_WDATA,
  SLAVE14_WSTRB,
  SLAVE14_WLAST,
  SLAVE14_WUSER,
  SLAVE14_WVALID,
  SLAVE14_WREADY,  

  SLAVE15_WID,
  SLAVE15_WDATA,
  SLAVE15_WSTRB,
  SLAVE15_WLAST,
  SLAVE15_WUSER,
  SLAVE15_WVALID,
  SLAVE15_WREADY,  

  SLAVE16_WID,
  SLAVE16_WDATA,
  SLAVE16_WSTRB,
  SLAVE16_WLAST,
  SLAVE16_WUSER,
  SLAVE16_WVALID,
  SLAVE16_WREADY,  

  SLAVE17_WID,
  SLAVE17_WDATA,
  SLAVE17_WSTRB,
  SLAVE17_WLAST,
  SLAVE17_WUSER,
  SLAVE17_WVALID,
  SLAVE17_WREADY,  

  SLAVE18_WID,
  SLAVE18_WDATA,
  SLAVE18_WSTRB,
  SLAVE18_WLAST,
  SLAVE18_WUSER,
  SLAVE18_WVALID,
  SLAVE18_WREADY,  

  SLAVE19_WID,
  SLAVE19_WDATA,
  SLAVE19_WSTRB,
  SLAVE19_WLAST,
  SLAVE19_WUSER,
  SLAVE19_WVALID,
  SLAVE19_WREADY,  

  SLAVE20_WID,
  SLAVE20_WDATA,
  SLAVE20_WSTRB,
  SLAVE20_WLAST,
  SLAVE20_WUSER,
  SLAVE20_WVALID,
  SLAVE20_WREADY,  

  SLAVE21_WID,
  SLAVE21_WDATA,
  SLAVE21_WSTRB,
  SLAVE21_WLAST,
  SLAVE21_WUSER,
  SLAVE21_WVALID,
  SLAVE21_WREADY,  

  SLAVE22_WID,
  SLAVE22_WDATA,
  SLAVE22_WSTRB,
  SLAVE22_WLAST,
  SLAVE22_WUSER,
  SLAVE22_WVALID,
  SLAVE22_WREADY,  

  SLAVE23_WID,
  SLAVE23_WDATA,
  SLAVE23_WSTRB,
  SLAVE23_WLAST,
  SLAVE23_WUSER,
  SLAVE23_WVALID,
  SLAVE23_WREADY,  

  SLAVE24_WID,
  SLAVE24_WDATA,
  SLAVE24_WSTRB,
  SLAVE24_WLAST,
  SLAVE24_WUSER,
  SLAVE24_WVALID,
  SLAVE24_WREADY,  

  SLAVE25_WID,
  SLAVE25_WDATA,
  SLAVE25_WSTRB,
  SLAVE25_WLAST,
  SLAVE25_WUSER,
  SLAVE25_WVALID,
  SLAVE25_WREADY,  

  SLAVE26_WID,
  SLAVE26_WDATA,
  SLAVE26_WSTRB,
  SLAVE26_WLAST,
  SLAVE26_WUSER,
  SLAVE26_WVALID,
  SLAVE26_WREADY,  

  SLAVE27_WID,
  SLAVE27_WDATA,
  SLAVE27_WSTRB,
  SLAVE27_WLAST,
  SLAVE27_WUSER,
  SLAVE27_WVALID,
  SLAVE27_WREADY,  

  SLAVE28_WID,
  SLAVE28_WDATA,
  SLAVE28_WSTRB,
  SLAVE28_WLAST,
  SLAVE28_WUSER,
  SLAVE28_WVALID,
  SLAVE28_WREADY,  

  SLAVE29_WID,
  SLAVE29_WDATA,
  SLAVE29_WSTRB,
  SLAVE29_WLAST,
  SLAVE29_WUSER,
  SLAVE29_WVALID,
  SLAVE29_WREADY,  

  SLAVE30_WID,
  SLAVE30_WDATA,
  SLAVE30_WSTRB,
  SLAVE30_WLAST,
  SLAVE30_WUSER,
  SLAVE30_WVALID,
  SLAVE30_WREADY,  

  SLAVE31_WID,
  SLAVE31_WDATA,
  SLAVE31_WSTRB,
  SLAVE31_WLAST,
  SLAVE31_WUSER,
  SLAVE31_WVALID,
  SLAVE31_WREADY,  
  
  // Slave Write Response Ports
  SLAVE0_BID,
  SLAVE0_BRESP,
  SLAVE0_BUSER,
  SLAVE0_BVALID,
  SLAVE0_BREADY,
   
   SLAVE1_BID,
  SLAVE1_BRESP,
  SLAVE1_BUSER,
  SLAVE1_BVALID,
  SLAVE1_BREADY,  
   
  SLAVE2_BID,
  SLAVE2_BRESP,
  SLAVE2_BUSER,
  SLAVE2_BVALID,
  SLAVE2_BREADY,
   
  SLAVE3_BID,
  SLAVE3_BRESP,
  SLAVE3_BUSER,
  SLAVE3_BVALID,
  SLAVE3_BREADY,
   
   SLAVE4_BID,
  SLAVE4_BRESP,
  SLAVE4_BUSER,
  SLAVE4_BVALID,
  SLAVE4_BREADY,  
   
   SLAVE5_BID,
  SLAVE5_BRESP,
  SLAVE5_BUSER,
  SLAVE5_BVALID,
  SLAVE5_BREADY,  
 
  SLAVE6_BID,
  SLAVE6_BRESP,
  SLAVE6_BUSER,
  SLAVE6_BVALID,
  SLAVE6_BREADY, 
 
  SLAVE7_BID,
  SLAVE7_BRESP,
  SLAVE7_BUSER,
  SLAVE7_BVALID,
  SLAVE7_BREADY,  
 
  SLAVE8_BID,
  SLAVE8_BRESP,
  SLAVE8_BUSER,
  SLAVE8_BVALID,
  SLAVE8_BREADY,  
 
  SLAVE9_BID,
  SLAVE9_BRESP,
  SLAVE9_BUSER,
  SLAVE9_BVALID,
  SLAVE9_BREADY,  
 
  SLAVE10_BID,
  SLAVE10_BRESP,
  SLAVE10_BUSER,
  SLAVE10_BVALID,
  SLAVE10_BREADY,  
 
  SLAVE11_BID,
  SLAVE11_BRESP,
  SLAVE11_BUSER,
  SLAVE11_BVALID,
  SLAVE11_BREADY,  
 
  SLAVE12_BID,
  SLAVE12_BRESP,
  SLAVE12_BUSER,
  SLAVE12_BVALID,
  SLAVE12_BREADY,  
 
  SLAVE13_BID,
  SLAVE13_BRESP,
  SLAVE13_BUSER,
  SLAVE13_BVALID,
  SLAVE13_BREADY,  
 
  SLAVE14_BID,
  SLAVE14_BRESP,
  SLAVE14_BUSER,
  SLAVE14_BVALID,
  SLAVE14_BREADY,  
 
  SLAVE15_BID,
  SLAVE15_BRESP,
  SLAVE15_BUSER,
  SLAVE15_BVALID,
  SLAVE15_BREADY,  
 
  SLAVE16_BID,
  SLAVE16_BRESP,
  SLAVE16_BUSER,
  SLAVE16_BVALID,
  SLAVE16_BREADY,  
 
  SLAVE17_BID,
  SLAVE17_BRESP,
  SLAVE17_BUSER,
  SLAVE17_BVALID,
  SLAVE17_BREADY,  
 
  SLAVE18_BID,
  SLAVE18_BRESP,
  SLAVE18_BUSER,
  SLAVE18_BVALID,
  SLAVE18_BREADY,  
 
  SLAVE19_BID,
  SLAVE19_BRESP,
  SLAVE19_BUSER,
  SLAVE19_BVALID,
  SLAVE19_BREADY,  
 
  SLAVE20_BID,
  SLAVE20_BRESP,
  SLAVE20_BUSER,
  SLAVE20_BVALID,
  SLAVE20_BREADY,  
 
  SLAVE21_BID,
  SLAVE21_BRESP,
  SLAVE21_BUSER,
  SLAVE21_BVALID,
  SLAVE21_BREADY,  
 
  SLAVE22_BID,
  SLAVE22_BRESP,
  SLAVE22_BUSER,
  SLAVE22_BVALID,
  SLAVE22_BREADY,  
 
  SLAVE23_BID,
  SLAVE23_BRESP,
  SLAVE23_BUSER,
  SLAVE23_BVALID,
  SLAVE23_BREADY,  
 
  SLAVE24_BID,
  SLAVE24_BRESP,
  SLAVE24_BUSER,
  SLAVE24_BVALID,
  SLAVE24_BREADY,  
 
  SLAVE25_BID,
  SLAVE25_BRESP,
  SLAVE25_BUSER,
  SLAVE25_BVALID,
  SLAVE25_BREADY,  
 
  SLAVE26_BID,
  SLAVE26_BRESP,
  SLAVE26_BUSER,
  SLAVE26_BVALID,
  SLAVE26_BREADY,   
 
  SLAVE27_BID,
  SLAVE27_BRESP,
  SLAVE27_BUSER,
  SLAVE27_BVALID,
  SLAVE27_BREADY,   
 
  SLAVE28_BID,
  SLAVE28_BRESP,
  SLAVE28_BUSER,
  SLAVE28_BVALID,
  SLAVE28_BREADY,   
 
  SLAVE29_BID,
  SLAVE29_BRESP,
  SLAVE29_BUSER,
  SLAVE29_BVALID,
  SLAVE29_BREADY,   
 
  SLAVE30_BID,
  SLAVE30_BRESP,
  SLAVE30_BUSER,
  SLAVE30_BVALID,
  SLAVE30_BREADY,   
 
  SLAVE31_BID,
  SLAVE31_BRESP,
  SLAVE31_BUSER,
  SLAVE31_BVALID,
  SLAVE31_BREADY, 
   
   // Slave Read Address Port
  SLAVE0_ARID,
  SLAVE0_ARADDR,
  SLAVE0_ARLEN,
  SLAVE0_ARSIZE,
  SLAVE0_ARBURST,
  SLAVE0_ARLOCK,
  SLAVE0_ARCACHE,
  SLAVE0_ARPROT,
  SLAVE0_ARREGION,    // not used
  SLAVE0_ARQOS,      // not used
  SLAVE0_ARUSER,
  SLAVE0_ARVALID,
  SLAVE0_ARREADY,
 
  SLAVE1_ARID,
  SLAVE1_ARADDR,
  SLAVE1_ARLEN,
  SLAVE1_ARSIZE,
  SLAVE1_ARBURST,
  SLAVE1_ARLOCK,
  SLAVE1_ARCACHE,
  SLAVE1_ARPROT,
  SLAVE1_ARREGION,    // not used
  SLAVE1_ARQOS,      // not used
  SLAVE1_ARUSER,
  SLAVE1_ARVALID,
  SLAVE1_ARREADY,

  SLAVE2_ARID,
  SLAVE2_ARADDR,
  SLAVE2_ARLEN,
  SLAVE2_ARSIZE,
  SLAVE2_ARBURST,
  SLAVE2_ARLOCK,
  SLAVE2_ARCACHE,
  SLAVE2_ARPROT,
  SLAVE2_ARREGION,    // not used
  SLAVE2_ARQOS,      // not used
  SLAVE2_ARUSER,
  SLAVE2_ARVALID,
  SLAVE2_ARREADY,

  SLAVE3_ARID,
  SLAVE3_ARADDR,
  SLAVE3_ARLEN,
  SLAVE3_ARSIZE,
  SLAVE3_ARBURST,
  SLAVE3_ARLOCK,
  SLAVE3_ARCACHE,
  SLAVE3_ARPROT,
  SLAVE3_ARREGION,    // not used
  SLAVE3_ARQOS,      // not used
  SLAVE3_ARUSER,
  SLAVE3_ARVALID,
  SLAVE3_ARREADY,

  SLAVE4_ARID,
  SLAVE4_ARADDR,
  SLAVE4_ARLEN,
  SLAVE4_ARSIZE,
  SLAVE4_ARBURST,
  SLAVE4_ARLOCK,
  SLAVE4_ARCACHE,
  SLAVE4_ARPROT,
  SLAVE4_ARREGION,    // not used
  SLAVE4_ARQOS,      // not used
  SLAVE4_ARUSER,
  SLAVE4_ARVALID,
  SLAVE4_ARREADY,

  SLAVE5_ARID,
  SLAVE5_ARADDR,
  SLAVE5_ARLEN,
  SLAVE5_ARSIZE,
  SLAVE5_ARBURST,
  SLAVE5_ARLOCK,
  SLAVE5_ARCACHE,
  SLAVE5_ARPROT,
  SLAVE5_ARREGION,    // not used
  SLAVE5_ARQOS,      // not used
  SLAVE5_ARUSER,
  SLAVE5_ARVALID,
  SLAVE5_ARREADY,
  
  SLAVE6_ARID,
  SLAVE6_ARADDR,
  SLAVE6_ARLEN,
  SLAVE6_ARSIZE,
  SLAVE6_ARBURST,
  SLAVE6_ARLOCK,
  SLAVE6_ARCACHE,
  SLAVE6_ARPROT,
  SLAVE6_ARREGION,    // not used
  SLAVE6_ARQOS,      // not used
  SLAVE6_ARUSER,
  SLAVE6_ARVALID,
  SLAVE6_ARREADY,  
  
  SLAVE7_ARID,
  SLAVE7_ARADDR,
  SLAVE7_ARLEN,
  SLAVE7_ARSIZE,
  SLAVE7_ARBURST,
  SLAVE7_ARLOCK,
  SLAVE7_ARCACHE,
  SLAVE7_ARPROT,
  SLAVE7_ARREGION,    // not used
  SLAVE7_ARQOS,      // not used
  SLAVE7_ARUSER,
  SLAVE7_ARVALID,
  SLAVE7_ARREADY,  
  
  SLAVE8_ARID,
  SLAVE8_ARADDR,
  SLAVE8_ARLEN,
  SLAVE8_ARSIZE,
  SLAVE8_ARBURST,
  SLAVE8_ARLOCK,
  SLAVE8_ARCACHE,
  SLAVE8_ARPROT,
  SLAVE8_ARREGION,    // not used
  SLAVE8_ARQOS,      // not used
  SLAVE8_ARUSER,
  SLAVE8_ARVALID,
  SLAVE8_ARREADY,  
  
  SLAVE9_ARID,
  SLAVE9_ARADDR,
  SLAVE9_ARLEN,
  SLAVE9_ARSIZE,
  SLAVE9_ARBURST,
  SLAVE9_ARLOCK,
  SLAVE9_ARCACHE,
  SLAVE9_ARPROT,
  SLAVE9_ARREGION,    // not used
  SLAVE9_ARQOS,      // not used
  SLAVE9_ARUSER,
  SLAVE9_ARVALID,
  SLAVE9_ARREADY,  
  
  SLAVE10_ARID,
  SLAVE10_ARADDR,
  SLAVE10_ARLEN,
  SLAVE10_ARSIZE,
  SLAVE10_ARBURST,
  SLAVE10_ARLOCK,
  SLAVE10_ARCACHE,
  SLAVE10_ARPROT,
  SLAVE10_ARREGION,    // not used
  SLAVE10_ARQOS,      // not used
  SLAVE10_ARUSER,
  SLAVE10_ARVALID,
  SLAVE10_ARREADY,  
  
  SLAVE11_ARID,
  SLAVE11_ARADDR,
  SLAVE11_ARLEN,
  SLAVE11_ARSIZE,
  SLAVE11_ARBURST,
  SLAVE11_ARLOCK,
  SLAVE11_ARCACHE,
  SLAVE11_ARPROT,
  SLAVE11_ARREGION,    // not used
  SLAVE11_ARQOS,      // not used
  SLAVE11_ARUSER,
  SLAVE11_ARVALID,
  SLAVE11_ARREADY,  
  
  SLAVE12_ARID,
  SLAVE12_ARADDR,
  SLAVE12_ARLEN,
  SLAVE12_ARSIZE,
  SLAVE12_ARBURST,
  SLAVE12_ARLOCK,
  SLAVE12_ARCACHE,
  SLAVE12_ARPROT,
  SLAVE12_ARREGION,    // not used
  SLAVE12_ARQOS,      // not used
  SLAVE12_ARUSER,
  SLAVE12_ARVALID,
  SLAVE12_ARREADY,  
  
  SLAVE13_ARID,
  SLAVE13_ARADDR,
  SLAVE13_ARLEN,
  SLAVE13_ARSIZE,
  SLAVE13_ARBURST,
  SLAVE13_ARLOCK,
  SLAVE13_ARCACHE,
  SLAVE13_ARPROT,
  SLAVE13_ARREGION,    // not used
  SLAVE13_ARQOS,      // not used
  SLAVE13_ARUSER,
  SLAVE13_ARVALID,
  SLAVE13_ARREADY,  
  
  SLAVE14_ARID,
  SLAVE14_ARADDR,
  SLAVE14_ARLEN,
  SLAVE14_ARSIZE,
  SLAVE14_ARBURST,
  SLAVE14_ARLOCK,
  SLAVE14_ARCACHE,
  SLAVE14_ARPROT,
  SLAVE14_ARREGION,    // not used
  SLAVE14_ARQOS,      // not used
  SLAVE14_ARUSER,
  SLAVE14_ARVALID,
  SLAVE14_ARREADY,  
  
  SLAVE15_ARID,
  SLAVE15_ARADDR,
  SLAVE15_ARLEN,
  SLAVE15_ARSIZE,
  SLAVE15_ARBURST,
  SLAVE15_ARLOCK,
  SLAVE15_ARCACHE,
  SLAVE15_ARPROT,
  SLAVE15_ARREGION,    // not used
  SLAVE15_ARQOS,      // not used
  SLAVE15_ARUSER,
  SLAVE15_ARVALID,
  SLAVE15_ARREADY,  
  
  SLAVE16_ARID,
  SLAVE16_ARADDR,
  SLAVE16_ARLEN,
  SLAVE16_ARSIZE,
  SLAVE16_ARBURST,
  SLAVE16_ARLOCK,
  SLAVE16_ARCACHE,
  SLAVE16_ARPROT,
  SLAVE16_ARREGION,    // not used
  SLAVE16_ARQOS,      // not used
  SLAVE16_ARUSER,
  SLAVE16_ARVALID,
  SLAVE16_ARREADY,  
  
  SLAVE17_ARID,
  SLAVE17_ARADDR,
  SLAVE17_ARLEN,
  SLAVE17_ARSIZE,
  SLAVE17_ARBURST,
  SLAVE17_ARLOCK,
  SLAVE17_ARCACHE,
  SLAVE17_ARPROT,
  SLAVE17_ARREGION,    // not used
  SLAVE17_ARQOS,      // not used
  SLAVE17_ARUSER,
  SLAVE17_ARVALID,
  SLAVE17_ARREADY,  
  
  SLAVE18_ARID,
  SLAVE18_ARADDR,
  SLAVE18_ARLEN,
  SLAVE18_ARSIZE,
  SLAVE18_ARBURST,
  SLAVE18_ARLOCK,
  SLAVE18_ARCACHE,
  SLAVE18_ARPROT,
  SLAVE18_ARREGION,    // not used
  SLAVE18_ARQOS,      // not used
  SLAVE18_ARUSER,
  SLAVE18_ARVALID,
  SLAVE18_ARREADY,  
  
  SLAVE19_ARID,
  SLAVE19_ARADDR,
  SLAVE19_ARLEN,
  SLAVE19_ARSIZE,
  SLAVE19_ARBURST,
  SLAVE19_ARLOCK,
  SLAVE19_ARCACHE,
  SLAVE19_ARPROT,
  SLAVE19_ARREGION,    // not used
  SLAVE19_ARQOS,      // not used
  SLAVE19_ARUSER,
  SLAVE19_ARVALID,
  SLAVE19_ARREADY,  
  
  SLAVE20_ARID,
  SLAVE20_ARADDR,
  SLAVE20_ARLEN,
  SLAVE20_ARSIZE,
  SLAVE20_ARBURST,
  SLAVE20_ARLOCK,
  SLAVE20_ARCACHE,
  SLAVE20_ARPROT,
  SLAVE20_ARREGION,    // not used
  SLAVE20_ARQOS,      // not used
  SLAVE20_ARUSER,
  SLAVE20_ARVALID,
  SLAVE20_ARREADY,  
  
  SLAVE21_ARID,
  SLAVE21_ARADDR,
  SLAVE21_ARLEN,
  SLAVE21_ARSIZE,
  SLAVE21_ARBURST,
  SLAVE21_ARLOCK,
  SLAVE21_ARCACHE,
  SLAVE21_ARPROT,
  SLAVE21_ARREGION,    // not used
  SLAVE21_ARQOS,      // not used
  SLAVE21_ARUSER,
  SLAVE21_ARVALID,
  SLAVE21_ARREADY,  
  
  SLAVE22_ARID,
  SLAVE22_ARADDR,
  SLAVE22_ARLEN,
  SLAVE22_ARSIZE,
  SLAVE22_ARBURST,
  SLAVE22_ARLOCK,
  SLAVE22_ARCACHE,
  SLAVE22_ARPROT,
  SLAVE22_ARREGION,    // not used
  SLAVE22_ARQOS,      // not used
  SLAVE22_ARUSER,
  SLAVE22_ARVALID,
  SLAVE22_ARREADY,    
  
  SLAVE23_ARID,
  SLAVE23_ARADDR,
  SLAVE23_ARLEN,
  SLAVE23_ARSIZE,
  SLAVE23_ARBURST,
  SLAVE23_ARLOCK,
  SLAVE23_ARCACHE,
  SLAVE23_ARPROT,
  SLAVE23_ARREGION,    // not used
  SLAVE23_ARQOS,      // not used
  SLAVE23_ARUSER,
  SLAVE23_ARVALID,
  SLAVE23_ARREADY,    
  
  SLAVE24_ARID,
  SLAVE24_ARADDR,
  SLAVE24_ARLEN,
  SLAVE24_ARSIZE,
  SLAVE24_ARBURST,
  SLAVE24_ARLOCK,
  SLAVE24_ARCACHE,
  SLAVE24_ARPROT,
  SLAVE24_ARREGION,    // not used
  SLAVE24_ARQOS,      // not used
  SLAVE24_ARUSER,
  SLAVE24_ARVALID,
  SLAVE24_ARREADY,    
  
  SLAVE25_ARID,
  SLAVE25_ARADDR,
  SLAVE25_ARLEN,
  SLAVE25_ARSIZE,
  SLAVE25_ARBURST,
  SLAVE25_ARLOCK,
  SLAVE25_ARCACHE,
  SLAVE25_ARPROT,
  SLAVE25_ARREGION,    // not used
  SLAVE25_ARQOS,      // not used
  SLAVE25_ARUSER,
  SLAVE25_ARVALID,
  SLAVE25_ARREADY,    
  
  SLAVE26_ARID,
  SLAVE26_ARADDR,
  SLAVE26_ARLEN,
  SLAVE26_ARSIZE,
  SLAVE26_ARBURST,
  SLAVE26_ARLOCK,
  SLAVE26_ARCACHE,
  SLAVE26_ARPROT,
  SLAVE26_ARREGION,    // not used
  SLAVE26_ARQOS,      // not used
  SLAVE26_ARUSER,
  SLAVE26_ARVALID,
  SLAVE26_ARREADY,    
  
  SLAVE27_ARID,
  SLAVE27_ARADDR,
  SLAVE27_ARLEN,
  SLAVE27_ARSIZE,
  SLAVE27_ARBURST,
  SLAVE27_ARLOCK,
  SLAVE27_ARCACHE,
  SLAVE27_ARPROT,
  SLAVE27_ARREGION,    // not used
  SLAVE27_ARQOS,      // not used
  SLAVE27_ARUSER,
  SLAVE27_ARVALID,
  SLAVE27_ARREADY,    
  
  SLAVE28_ARID,
  SLAVE28_ARADDR,
  SLAVE28_ARLEN,
  SLAVE28_ARSIZE,
  SLAVE28_ARBURST,
  SLAVE28_ARLOCK,
  SLAVE28_ARCACHE,
  SLAVE28_ARPROT,
  SLAVE28_ARREGION,    // not used
  SLAVE28_ARQOS,      // not used
  SLAVE28_ARUSER,
  SLAVE28_ARVALID,
  SLAVE28_ARREADY,    
  
  SLAVE29_ARID,
  SLAVE29_ARADDR,
  SLAVE29_ARLEN,
  SLAVE29_ARSIZE,
  SLAVE29_ARBURST,
  SLAVE29_ARLOCK,
  SLAVE29_ARCACHE,
  SLAVE29_ARPROT,
  SLAVE29_ARREGION,    // not used
  SLAVE29_ARQOS,      // not used
  SLAVE29_ARUSER,
  SLAVE29_ARVALID,
  SLAVE29_ARREADY,    
  
  SLAVE30_ARID,
  SLAVE30_ARADDR,
  SLAVE30_ARLEN,
  SLAVE30_ARSIZE,
  SLAVE30_ARBURST,
  SLAVE30_ARLOCK,
  SLAVE30_ARCACHE,
  SLAVE30_ARPROT,
  SLAVE30_ARREGION,    // not used
  SLAVE30_ARQOS,      // not used
  SLAVE30_ARUSER,
  SLAVE30_ARVALID,
  SLAVE30_ARREADY,    
  
  SLAVE31_ARID,
  SLAVE31_ARADDR,
  SLAVE31_ARLEN,
  SLAVE31_ARSIZE,
  SLAVE31_ARBURST,
  SLAVE31_ARLOCK,
  SLAVE31_ARCACHE,
  SLAVE31_ARPROT,
  SLAVE31_ARREGION,    // not used
  SLAVE31_ARQOS,      // not used
  SLAVE31_ARUSER,
  SLAVE31_ARVALID,
  SLAVE31_ARREADY,  
  
   // Slave Read Data Ports
  SLAVE0_RID,
  SLAVE0_RDATA,
  SLAVE0_RRESP,
  SLAVE0_RLAST,
  SLAVE0_RUSER,      // not used
  SLAVE0_RVALID,
  SLAVE0_RREADY,
   
  SLAVE1_RID,
  SLAVE1_RDATA,
  SLAVE1_RRESP,
  SLAVE1_RLAST,
  SLAVE1_RUSER,      // not used
  SLAVE1_RVALID,
  SLAVE1_RREADY,   
   
  SLAVE2_RID,
  SLAVE2_RDATA,
  SLAVE2_RRESP,
  SLAVE2_RLAST,
  SLAVE2_RUSER,      // not used
  SLAVE2_RVALID,
  SLAVE2_RREADY,   
 
  SLAVE3_RID,
  SLAVE3_RDATA,
  SLAVE3_RRESP,
  SLAVE3_RLAST,
  SLAVE3_RUSER,      // not used
  SLAVE3_RVALID,
  SLAVE3_RREADY, 
   
  SLAVE4_RID,
  SLAVE4_RDATA,
  SLAVE4_RRESP,
  SLAVE4_RLAST,
  SLAVE4_RUSER,      // not used
  SLAVE4_RVALID,
  SLAVE4_RREADY,   
   
  SLAVE5_RID,
  SLAVE5_RDATA,
  SLAVE5_RRESP,
  SLAVE5_RLAST,
  SLAVE5_RUSER,      // not used
  SLAVE5_RVALID,
  SLAVE5_RREADY,   
   
  SLAVE6_RID,
  SLAVE6_RDATA,
  SLAVE6_RRESP,
  SLAVE6_RLAST,
  SLAVE6_RUSER,      // not used
  SLAVE6_RVALID,
  SLAVE6_RREADY,
   
  SLAVE7_RID,
  SLAVE7_RDATA,
  SLAVE7_RRESP,
  SLAVE7_RLAST,
  SLAVE7_RUSER,      // not used
  SLAVE7_RVALID,
  SLAVE7_RREADY,
   
  SLAVE8_RID,
  SLAVE8_RDATA,
  SLAVE8_RRESP,
  SLAVE8_RLAST,
  SLAVE8_RUSER,      // not used
  SLAVE8_RVALID,
  SLAVE8_RREADY,
   
  SLAVE9_RID,
  SLAVE9_RDATA,
  SLAVE9_RRESP,
  SLAVE9_RLAST,
  SLAVE9_RUSER,      // not used
  SLAVE9_RVALID,
  SLAVE9_RREADY,
   
  SLAVE10_RID,
  SLAVE10_RDATA,
  SLAVE10_RRESP,
  SLAVE10_RLAST,
  SLAVE10_RUSER,      // not used
  SLAVE10_RVALID,
  SLAVE10_RREADY,
   
  SLAVE11_RID,
  SLAVE11_RDATA,
  SLAVE11_RRESP,
  SLAVE11_RLAST,
  SLAVE11_RUSER,      // not used
  SLAVE11_RVALID,
  SLAVE11_RREADY,
   
  SLAVE12_RID,
  SLAVE12_RDATA,
  SLAVE12_RRESP,
  SLAVE12_RLAST,
  SLAVE12_RUSER,      // not used
  SLAVE12_RVALID,
  SLAVE12_RREADY,
   
  SLAVE13_RID,
  SLAVE13_RDATA,
  SLAVE13_RRESP,
  SLAVE13_RLAST,
  SLAVE13_RUSER,      // not used
  SLAVE13_RVALID,
  SLAVE13_RREADY,
   
  SLAVE14_RID,
  SLAVE14_RDATA,
  SLAVE14_RRESP,
  SLAVE14_RLAST,
  SLAVE14_RUSER,      // not used
  SLAVE14_RVALID,
  SLAVE14_RREADY,
   
  SLAVE15_RID,
  SLAVE15_RDATA,
  SLAVE15_RRESP,
  SLAVE15_RLAST,
  SLAVE15_RUSER,      // not used
  SLAVE15_RVALID,
  SLAVE15_RREADY,
   
  SLAVE16_RID,
  SLAVE16_RDATA,
  SLAVE16_RRESP,
  SLAVE16_RLAST,
  SLAVE16_RUSER,      // not used
  SLAVE16_RVALID,
  SLAVE16_RREADY,
   
  SLAVE17_RID,
  SLAVE17_RDATA,
  SLAVE17_RRESP,
  SLAVE17_RLAST,
  SLAVE17_RUSER,      // not used
  SLAVE17_RVALID,
  SLAVE17_RREADY,
   
  SLAVE18_RID,
  SLAVE18_RDATA,
  SLAVE18_RRESP,
  SLAVE18_RLAST,
  SLAVE18_RUSER,      // not used
  SLAVE18_RVALID,
  SLAVE18_RREADY,
   
  SLAVE19_RID,
  SLAVE19_RDATA,
  SLAVE19_RRESP,
  SLAVE19_RLAST,
  SLAVE19_RUSER,      // not used
  SLAVE19_RVALID,
  SLAVE19_RREADY,
   
  SLAVE20_RID,
  SLAVE20_RDATA,
  SLAVE20_RRESP,
  SLAVE20_RLAST,
  SLAVE20_RUSER,      // not used
  SLAVE20_RVALID,
  SLAVE20_RREADY,
   
  SLAVE21_RID,
  SLAVE21_RDATA,
  SLAVE21_RRESP,
  SLAVE21_RLAST,
  SLAVE21_RUSER,      // not used
  SLAVE21_RVALID,
  SLAVE21_RREADY,
   
  SLAVE22_RID,
  SLAVE22_RDATA,
  SLAVE22_RRESP,
  SLAVE22_RLAST,
  SLAVE22_RUSER,      // not used
  SLAVE22_RVALID,
  SLAVE22_RREADY,
   
  SLAVE23_RID,
  SLAVE23_RDATA,
  SLAVE23_RRESP,
  SLAVE23_RLAST,
  SLAVE23_RUSER,      // not used
  SLAVE23_RVALID,
  SLAVE23_RREADY,
   
  SLAVE24_RID,
  SLAVE24_RDATA,
  SLAVE24_RRESP,
  SLAVE24_RLAST,
  SLAVE24_RUSER,      // not used
  SLAVE24_RVALID,
  SLAVE24_RREADY,
   
  SLAVE25_RID,
  SLAVE25_RDATA,
  SLAVE25_RRESP,
  SLAVE25_RLAST,
  SLAVE25_RUSER,      // not used
  SLAVE25_RVALID,
  SLAVE25_RREADY,
   
  SLAVE26_RID,
  SLAVE26_RDATA,
  SLAVE26_RRESP,
  SLAVE26_RLAST,
  SLAVE26_RUSER,      // not used
  SLAVE26_RVALID,
  SLAVE26_RREADY,
   
  SLAVE27_RID,
  SLAVE27_RDATA,
  SLAVE27_RRESP,
  SLAVE27_RLAST,
  SLAVE27_RUSER,      // not used
  SLAVE27_RVALID,
  SLAVE27_RREADY,
   
  SLAVE28_RID,
  SLAVE28_RDATA,
  SLAVE28_RRESP,
  SLAVE28_RLAST,
  SLAVE28_RUSER,      // not used
  SLAVE28_RVALID,
  SLAVE28_RREADY,
   
  SLAVE29_RID,
  SLAVE29_RDATA,
  SLAVE29_RRESP,
  SLAVE29_RLAST,
  SLAVE29_RUSER,      // not used
  SLAVE29_RVALID,
  SLAVE29_RREADY,
   
  SLAVE30_RID,
  SLAVE30_RDATA,
  SLAVE30_RRESP,
  SLAVE30_RLAST,
  SLAVE30_RUSER,      // not used
  SLAVE30_RVALID,
  SLAVE30_RREADY,
   
  SLAVE31_RID,
  SLAVE31_RDATA,
  SLAVE31_RRESP,
  SLAVE31_RLAST,
  SLAVE31_RUSER,      // not used
  SLAVE31_RVALID,
  SLAVE31_RREADY
  
   )
   
     /* jh_synthesis syn_hier = "flatten" */ ;
   
   //=====================================================================
   // Global Parameters
   //=====================================================================
   
  parameter integer FAMILY                = 19;
    
  parameter integer NUM_MASTERS      = 8;        // defines number of master ports 
  parameter integer NUM_SLAVES         = 8;        // defines number of slaves

  parameter integer ID_WIDTH         = 1;        // number of bits for ID (ie AID, WID, BID) - valid 1-8 
  parameter integer ADDR_WIDTH          = 20;        // valid values - 16 - 64

  //====================================================================
  // Crossbar parameters
  //====================================================================
  parameter integer DATA_WIDTH       = 32;        // valid widths - 32, 64, 128

  parameter NUM_THREADS          = 1;        // defined number of indpendent threads per master supported - valid range 1-8
  parameter OPEN_TRANS_MAX        = 2;        // max number of outstanding transactions per thread - valid range 1-8
    
  localparam OPEN_WRTRANS_MAX       = ($clog2(NUM_MASTERS*OPEN_TRANS_MAX*NUM_THREADS) > 2) ? $clog2(NUM_MASTERS*OPEN_TRANS_MAX*NUM_THREADS) : 2;        // max number of outstanding write transactions - valid range 2-8 - 2**OPEN_WRTRANS_MAX
  localparam OPEN_RDTRANS_MAX       = ($clog2(NUM_MASTERS*OPEN_TRANS_MAX*NUM_THREADS) > 2) ? $clog2(NUM_MASTERS*OPEN_TRANS_MAX*NUM_THREADS) : 2;        // max number of outstanding read transactions - valid range  2-8 - 2**OPEN_RDTRANS_MAX

  

/* 
  SAR 94407 Change Start  
  
  Below parameters are removed as a global parameters and used as a local parameter  
  
  parameter UPPER_COMPARE_BIT       = 15;        // Defines the upper bit of range to compare
  parameter LOWER_COMPARE_BIT       = 12;        // Defines lower bound of compare - bits below are dont care
  
  
  //Below parameters are removed as it is no longer used.As these parameters are used in RTL and to remove warnings/errors it is declared 
  //as local parameter 
 
  parameter [63:0]  SLOT0_BASE_VEC = 'h0;          // Defines the base address for Slave 0 decode
  parameter [63:0]  SLOT1_BASE_VEC = 'h1;          // Defines the base address for Slave 1 decode
  parameter [63:0]  SLOT2_BASE_VEC = 'h2;          // Defines the base address for Slave 2 decode
  parameter [63:0]  SLOT3_BASE_VEC = 'h3;          // Defines the base address for Slave 3 decode
  parameter [63:0]  SLOT4_BASE_VEC = 'h4;          // Defines the base address for Slave 4 decode
  parameter [63:0]  SLOT5_BASE_VEC = 'h5;          // Defines the base address for Slave 5 decode
  parameter [63:0]  SLOT6_BASE_VEC = 'h6;          // Defines the base address for Slave 6 decode
  parameter [63:0]  SLOT7_BASE_VEC = 'h7;          // Defines the base address for Slave 7 decode
  parameter [63:0]  SLOT8_BASE_VEC  = 'h8;          // Defines the base address for Slave 8 decode
  parameter [63:0]  SLOT9_BASE_VEC  = 'h9;          // Defines the base address for Slave 9 decode
  parameter [63:0]  SLOT10_BASE_VEC = 'ha;          // Defines the base address for Slave 10 decode
  parameter [63:0]  SLOT11_BASE_VEC = 'hb;          // Defines the base address for Slave 11 decode
  parameter [63:0]  SLOT12_BASE_VEC = 'hc;          // Defines the base address for Slave 12 decode
  parameter [63:0]  SLOT13_BASE_VEC = 'hd;          // Defines the base address for Slave 13 decode
  parameter [63:0]  SLOT14_BASE_VEC = 'he;          // Defines the base address for Slave 14 decode
  parameter [63:0]  SLOT15_BASE_VEC = 'hf;          // Defines the base address for Slave 15 decode
  parameter [63:0]  SLOT16_BASE_VEC = 'h10;          // Defines the base address for Slave 16 decode
  parameter [63:0]  SLOT17_BASE_VEC = 'h11;          // Defines the base address for Slave 17 decode
  parameter [63:0]  SLOT18_BASE_VEC = 'h12;          // Defines the base address for Slave 18 decode
  parameter [63:0]  SLOT19_BASE_VEC = 'h13;          // Defines the base address for Slave 19 decode
  parameter [63:0]  SLOT20_BASE_VEC = 'h14;          // Defines the base address for Slave 20 decode
  parameter [63:0]  SLOT21_BASE_VEC = 'h15;          // Defines the base address for Slave 21 decode
  parameter [63:0]  SLOT22_BASE_VEC = 'h16;          // Defines the base address for Slave 22 decode
  parameter [63:0]  SLOT23_BASE_VEC = 'h17;          // Defines the base address for Slave 23 decode
  parameter [63:0]  SLOT24_BASE_VEC = 'h18;          // Defines the base address for Slave 24 decode
  parameter [63:0]  SLOT25_BASE_VEC = 'h19;          // Defines the base address for Slave 25 decode
  parameter [63:0]  SLOT26_BASE_VEC = 'h1a;          // Defines the base address for Slave 26 decode
  parameter [63:0]  SLOT27_BASE_VEC = 'h1b;          // Defines the base address for Slave 27 decode
  parameter [63:0]  SLOT28_BASE_VEC = 'h1c;          // Defines the base address for Slave 28 decode
  parameter [63:0]  SLOT29_BASE_VEC = 'h1d;          // Defines the base address for Slave 29 decode
  parameter [63:0]  SLOT30_BASE_VEC = 'h1e;          // Defines the base address for Slave 30 decode
  parameter [63:0]  SLOT31_BASE_VEC = 'h1f;          // Defines the base address for Slave 31 decode

*/

  localparam [ADDR_WIDTH-1:0]  SLOT0_BASE_VEC = 'h0;          // Defines the base address for Slave 0 decode
  localparam [ADDR_WIDTH-1:0]  SLOT1_BASE_VEC = 'h1;          // Defines the base address for Slave 1 decode
  localparam [ADDR_WIDTH-1:0]  SLOT2_BASE_VEC = 'h2;          // Defines the base address for Slave 2 decode
  localparam [ADDR_WIDTH-1:0]  SLOT3_BASE_VEC = 'h3;          // Defines the base address for Slave 3 decode
  localparam [ADDR_WIDTH-1:0]  SLOT4_BASE_VEC = 'h4;          // Defines the base address for Slave 4 decode
  localparam [ADDR_WIDTH-1:0]  SLOT5_BASE_VEC = 'h5;          // Defines the base address for Slave 5 decode
  localparam [ADDR_WIDTH-1:0]  SLOT6_BASE_VEC = 'h6;          // Defines the base address for Slave 6 decode
  localparam [ADDR_WIDTH-1:0]  SLOT7_BASE_VEC = 'h7;          // Defines the base address for Slave 7 decode
  localparam [ADDR_WIDTH-1:0]  SLOT8_BASE_VEC  = 'h8;          // Defines the base address for Slave 8 decode
  localparam [ADDR_WIDTH-1:0]  SLOT9_BASE_VEC  = 'h9;          // Defines the base address for Slave 9 decode
  localparam [ADDR_WIDTH-1:0]  SLOT10_BASE_VEC = 'ha;          // Defines the base address for Slave 10 decode
  localparam [ADDR_WIDTH-1:0]  SLOT11_BASE_VEC = 'hb;          // Defines the base address for Slave 11 decode
  localparam [ADDR_WIDTH-1:0]  SLOT12_BASE_VEC = 'hc;          // Defines the base address for Slave 12 decode
  localparam [ADDR_WIDTH-1:0]  SLOT13_BASE_VEC = 'hd;          // Defines the base address for Slave 13 decode
  localparam [ADDR_WIDTH-1:0]  SLOT14_BASE_VEC = 'he;          // Defines the base address for Slave 14 decode
  localparam [ADDR_WIDTH-1:0]  SLOT15_BASE_VEC = 'hf;          // Defines the base address for Slave 15 decode
  localparam [ADDR_WIDTH-1:0]  SLOT16_BASE_VEC = 'h10;          // Defines the base address for Slave 16 decode
  localparam [ADDR_WIDTH-1:0]  SLOT17_BASE_VEC = 'h11;          // Defines the base address for Slave 17 decode
  localparam [ADDR_WIDTH-1:0]  SLOT18_BASE_VEC = 'h12;          // Defines the base address for Slave 18 decode
  localparam [ADDR_WIDTH-1:0]  SLOT19_BASE_VEC = 'h13;          // Defines the base address for Slave 19 decode
  localparam [ADDR_WIDTH-1:0]  SLOT20_BASE_VEC = 'h14;          // Defines the base address for Slave 20 decode
  localparam [ADDR_WIDTH-1:0]  SLOT21_BASE_VEC = 'h15;          // Defines the base address for Slave 21 decode
  localparam [ADDR_WIDTH-1:0]  SLOT22_BASE_VEC = 'h16;          // Defines the base address for Slave 22 decode
  localparam [ADDR_WIDTH-1:0]  SLOT23_BASE_VEC = 'h17;          // Defines the base address for Slave 23 decode
  localparam [ADDR_WIDTH-1:0]  SLOT24_BASE_VEC = 'h18;          // Defines the base address for Slave 24 decode
  localparam [ADDR_WIDTH-1:0]  SLOT25_BASE_VEC = 'h19;          // Defines the base address for Slave 25 decode
  localparam [ADDR_WIDTH-1:0]  SLOT26_BASE_VEC = 'h1a;          // Defines the base address for Slave 26 decode
  localparam [ADDR_WIDTH-1:0]  SLOT27_BASE_VEC = 'h1b;          // Defines the base address for Slave 27 decode
  localparam [ADDR_WIDTH-1:0]  SLOT28_BASE_VEC = 'h1c;          // Defines the base address for Slave 28 decode
  localparam [ADDR_WIDTH-1:0]  SLOT29_BASE_VEC = 'h1d;          // Defines the base address for Slave 29 decode
  localparam [ADDR_WIDTH-1:0]  SLOT30_BASE_VEC = 'h1e;          // Defines the base address for Slave 30 decode
  localparam [ADDR_WIDTH-1:0]  SLOT31_BASE_VEC = 'h1f;          // Defines the base address for Slave 31 decode
  
  //Following parameters used for MIN_VEC and MAX_VEC per slave are removed as a global parameters and used as a local parameters

/*  
  parameter [ADDR_WIDTH-1:0]   SLOT0_MIN_VEC  = 'h0;          // SLOT0 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT1_MIN_VEC  = 'h0;          // SLOT1 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT2_MIN_VEC  = 'h0;          // SLOT2 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT3_MIN_VEC  = 'h0;          // SLOT3 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT4_MIN_VEC  = 'h0;          // SLOT4 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT5_MIN_VEC  = 'h0;          // SLOT5 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT6_MIN_VEC  = 'h0;          // SLOT6 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT7_MIN_VEC  = 'h0;          // SLOT7 Min address
  parameter [ADDR_WIDTH-1:0]   SLOT8_MIN_VEC  = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT9_MIN_VEC  = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT10_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT11_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT12_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT13_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT14_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT15_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT16_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT17_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT18_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT19_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT20_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT21_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT22_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT23_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT24_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT25_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT26_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT27_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT28_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT29_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT30_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  parameter [ADDR_WIDTH-1:0]   SLOT31_MIN_VEC = 'h0;          // Defines the Min address for Slave 7 decode
  
  parameter [ADDR_WIDTH-1:0]   SLOT0_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT0 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT1_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT1 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT2_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT2 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT3_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT3 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT4_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT4 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT5_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT5 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT6_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT6 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT7_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT7 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT8_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT8 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT9_MAX_VEC  = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT9 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT10_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT10 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT11_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT11 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT12_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT12 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT13_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT13 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT14_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT14 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT15_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT15 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT16_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT16 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT17_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT17 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT18_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT18 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT19_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT19 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT20_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT20 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT21_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT21 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT22_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT22 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT23_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT23 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT24_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT24 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT25_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT25 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT26_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT26 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT27_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT27 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT28_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT28 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT29_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT29 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT30_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT30 Max address
  parameter [ADDR_WIDTH-1:0]   SLOT31_MAX_VEC = 64'hFFFF_FFFF_FFFF_FFFF;      // SLOT31 Max address
  
*/									     

  //SLOTy_START_ADDR parameter is added for each slave

  parameter [ADDR_WIDTH-1:0] SLAVE0_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE1_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE2_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE3_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE4_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE5_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE6_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE7_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE8_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE9_START_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE10_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE11_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE12_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE13_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE14_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE15_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE16_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE17_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE18_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE19_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE20_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE21_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE22_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE23_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE24_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE25_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE26_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE27_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE28_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE29_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE30_START_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE31_START_ADDR = {ADDR_WIDTH{1'b0}};

 //SLOTy_END_ADDR parameter is added for each slave 
  
  parameter [ADDR_WIDTH-1:0] SLAVE0_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE1_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE2_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE3_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE4_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE5_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE6_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE7_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE8_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE9_END_ADDR  = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE10_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE11_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE12_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE13_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE14_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE15_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE16_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE17_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE18_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE19_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE20_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE21_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE22_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE23_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE24_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE25_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE26_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE27_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE28_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE29_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE30_END_ADDR = {ADDR_WIDTH{1'b0}};
  parameter [ADDR_WIDTH-1:0] SLAVE31_END_ADDR = {ADDR_WIDTH{1'b0}};  

  //As new parameters SLAVE_START_ADDR and SLAVE_END_ADDR,UPPER_COMPARE_BIT and LOWER_COMPARE_BIT parameters are no longer required.
  //However to remove warnings/errors,UPPER_COMPARE_BIT is assigned to ADDR_WIDTH and LOWER_COMPARE_BIT is assigned to 0
  
  localparam UPPER_COMPARE_BIT = ADDR_WIDTH;
  localparam LOWER_COMPARE_BIT = 0;
  
  
  //Local parameter used to assign START ADDRESS for each slave to minimize the RTL Change
  
  localparam [ADDR_WIDTH-1: 0]   SLOT0_MIN_VEC  = SLAVE0_START_ADDR;           // SLOT0 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT1_MIN_VEC  = SLAVE1_START_ADDR;           // SLOT1 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT2_MIN_VEC  = SLAVE2_START_ADDR;           // SLOT2 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT3_MIN_VEC  = SLAVE3_START_ADDR;           // SLOT3 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT4_MIN_VEC  = SLAVE4_START_ADDR;           // SLOT4 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT5_MIN_VEC  = SLAVE5_START_ADDR;           // SLOT5 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT6_MIN_VEC  = SLAVE6_START_ADDR;           // SLOT6 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT7_MIN_VEC  = SLAVE7_START_ADDR;           // SLOT7 start address
  localparam [ADDR_WIDTH-1: 0]   SLOT8_MIN_VEC  = SLAVE8_START_ADDR;           // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT9_MIN_VEC  = SLAVE9_START_ADDR;           // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT10_MIN_VEC = SLAVE10_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT11_MIN_VEC = SLAVE11_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT12_MIN_VEC = SLAVE12_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT13_MIN_VEC = SLAVE13_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT14_MIN_VEC = SLAVE14_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT15_MIN_VEC = SLAVE15_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT16_MIN_VEC = SLAVE16_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT17_MIN_VEC = SLAVE17_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT18_MIN_VEC = SLAVE18_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT19_MIN_VEC = SLAVE19_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT20_MIN_VEC = SLAVE20_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT21_MIN_VEC = SLAVE21_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT22_MIN_VEC = SLAVE22_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT23_MIN_VEC = SLAVE23_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT24_MIN_VEC = SLAVE24_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT25_MIN_VEC = SLAVE25_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT26_MIN_VEC = SLAVE26_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT27_MIN_VEC = SLAVE27_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT28_MIN_VEC = SLAVE28_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT29_MIN_VEC = SLAVE29_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT30_MIN_VEC = SLAVE30_START_ADDR;          // Defines the start address for Slave 7 decode
  localparam [ADDR_WIDTH-1: 0]   SLOT31_MIN_VEC = SLAVE31_START_ADDR;          // Defines the start address for Slave 7 decode
  
  //Local parameter used to assign END ADDRESS for each slave to minimize the RTL Change
  
  localparam [ADDR_WIDTH-1: 0]   SLOT0_MAX_VEC  = SLAVE0_END_ADDR;           // SLOT0 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT1_MAX_VEC  = SLAVE1_END_ADDR;           // SLOT1 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT2_MAX_VEC  = SLAVE2_END_ADDR;           // SLOT2 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT3_MAX_VEC  = SLAVE3_END_ADDR;           // SLOT3 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT4_MAX_VEC  = SLAVE4_END_ADDR;           // SLOT4 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT5_MAX_VEC  = SLAVE5_END_ADDR;           // SLOT5 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT6_MAX_VEC  = SLAVE6_END_ADDR;           // SLOT6 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT7_MAX_VEC  = SLAVE7_END_ADDR;           // SLOT7 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT8_MAX_VEC  = SLAVE8_END_ADDR;           // SLOT8 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT9_MAX_VEC  = SLAVE9_END_ADDR;           // SLOT9 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT10_MAX_VEC = SLAVE10_END_ADDR;          // SLOT10 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT11_MAX_VEC = SLAVE11_END_ADDR;          // SLOT11 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT12_MAX_VEC = SLAVE12_END_ADDR;          // SLOT12 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT13_MAX_VEC = SLAVE13_END_ADDR;          // SLOT13 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT14_MAX_VEC = SLAVE14_END_ADDR;          // SLOT14 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT15_MAX_VEC = SLAVE15_END_ADDR;          // SLOT15 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT16_MAX_VEC = SLAVE16_END_ADDR;          // SLOT16 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT17_MAX_VEC = SLAVE17_END_ADDR;          // SLOT17 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT18_MAX_VEC = SLAVE18_END_ADDR;          // SLOT18 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT19_MAX_VEC = SLAVE19_END_ADDR;          // SLOT19 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT20_MAX_VEC = SLAVE20_END_ADDR;          // SLOT20 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT21_MAX_VEC = SLAVE21_END_ADDR;          // SLOT21 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT22_MAX_VEC = SLAVE22_END_ADDR;          // SLOT22 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT23_MAX_VEC = SLAVE23_END_ADDR;          // SLOT23 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT24_MAX_VEC = SLAVE24_END_ADDR;          // SLOT24 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT25_MAX_VEC = SLAVE25_END_ADDR;          // SLOT25 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT26_MAX_VEC = SLAVE26_END_ADDR;          // SLOT26 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT27_MAX_VEC = SLAVE27_END_ADDR;          // SLOT27 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT28_MAX_VEC = SLAVE28_END_ADDR;          // SLOT28 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT29_MAX_VEC = SLAVE29_END_ADDR;          // SLOT29 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT30_MAX_VEC = SLAVE30_END_ADDR;          // SLOT30 End address
  localparam [ADDR_WIDTH-1: 0]   SLOT31_MAX_VEC = SLAVE31_END_ADDR;          // SLOT31 End address
  
  //SAR 94407 Change End

  localparam integer SUPPORT_USER_SIGNALS   = 0;        // indicates where user signals upport - 0 mean no, 1 means yes
  parameter integer USER_WIDTH       = 1;               // defines the number of bits for USER signals RUSER and WUSER
  parameter integer CROSSBAR_MODE      = 1;             // defines whether non-blocking (ie set 1) or shared access data path

  parameter [0:0]    MASTER0_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port

  parameter [0:0]    MASTER0_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER0_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER0_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port
            
  parameter [0:0]    MASTER1_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port

  parameter [0:0]    MASTER1_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER1_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER1_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port

  parameter [0:0]    MASTER2_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port  

  parameter [0:0]    MASTER2_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER2_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER2_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port
            
  parameter [0:0]    MASTER3_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port  
  
  parameter [0:0]    MASTER3_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER3_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER3_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port
            
  parameter [0:0]    MASTER4_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port  

  parameter [0:0]    MASTER4_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER4_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER4_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port
            
  parameter [0:0]    MASTER5_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port  

  parameter [0:0]    MASTER5_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER5_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER5_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port
            
  parameter [0:0]    MASTER6_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port

  parameter [0:0]    MASTER6_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER6_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER6_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port
              
  parameter [0:0]    MASTER7_WRITE_SLAVE0  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE1  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE2  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE3  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE4  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE5  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE6  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE7  = 1'b1;      // bit for slave indicating if a master can write to that port

  parameter [0:0]    MASTER7_WRITE_SLAVE8  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE9  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE10  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE11  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE12  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE13  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE14  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE15  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE16  = 1'b1;      // bit for slave indicating if a master can write to that port  
  parameter [0:0]    MASTER7_WRITE_SLAVE17  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE18  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE19  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE20  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE21  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE22  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE23  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE24  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE25  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE26  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE27  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE28  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE29  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE30  = 1'b1;      // bit for slave indicating if a master can write to that port
  parameter [0:0]    MASTER7_WRITE_SLAVE31  = 1'b1;      // bit for slave indicating if a master can write to that port

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////              

  parameter [0:0]    MASTER0_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port

  parameter [0:0]    MASTER0_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER0_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER0_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port

  
  parameter [0:0]    MASTER1_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port

  parameter [0:0]    MASTER1_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER1_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER1_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port

  
  parameter [0:0]    MASTER2_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port  

  parameter [0:0]    MASTER2_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER2_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER2_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port     

  
  parameter [0:0]    MASTER3_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port  

  parameter [0:0]    MASTER3_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER3_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER3_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port 

  
  parameter [0:0]    MASTER4_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port  

  parameter [0:0]    MASTER4_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER4_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER4_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port 

  
  parameter [0:0]    MASTER5_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port  

  parameter [0:0]    MASTER5_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER5_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER5_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port 

  
  parameter [0:0]    MASTER6_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port

  parameter [0:0]    MASTER6_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER6_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER6_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port 

  
  parameter [0:0]    MASTER7_READ_SLAVE0  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE1  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE2  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE3  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE4  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE5  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE6  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE7  = 1'b1;      // bit for slave indicating if a master can read to that port

  parameter [0:0]    MASTER7_READ_SLAVE8  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE9  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE10  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE11  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE12  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE13  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE14  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE15  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE16  = 1'b1;      // bit for slave indicating if a master can read to that port  
  parameter [0:0]    MASTER7_READ_SLAVE17  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE18  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE19  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE20  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE21  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE22  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE23  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE24  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE25  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE26  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE27  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE28  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE29  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE30  = 1'b1;      // bit for slave indicating if a master can read to that port
  parameter [0:0]    MASTER7_READ_SLAVE31  = 1'b1;      // bit for slave indicating if a master can read to that port 

  parameter  RD_ARB_EN           = 1;        // select arb or ordered rdata

  parameter [0:0]  MASTER0_CLOCK_DOMAIN_CROSSING  = 1'b0;  
  parameter [0:0]  MASTER1_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  MASTER2_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  MASTER3_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  MASTER4_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  MASTER5_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  MASTER6_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  MASTER7_CLOCK_DOMAIN_CROSSING  = MASTER0_CLOCK_DOMAIN_CROSSING;    
  
  parameter [0:0]  SLAVE0_CLOCK_DOMAIN_CROSSING  = 1'b0;  
  parameter [0:0]  SLAVE1_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  SLAVE2_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  SLAVE3_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE4_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  SLAVE5_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  SLAVE6_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;  
  parameter [0:0]  SLAVE7_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;

  parameter [0:0]  SLAVE8_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE9_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE10_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE11_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE12_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE13_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE14_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE15_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE16_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE17_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE18_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE19_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE20_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE21_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE22_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE23_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE24_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE25_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE26_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE27_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE28_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE29_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE30_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;
  parameter [0:0]  SLAVE31_CLOCK_DOMAIN_CROSSING  = SLAVE0_CLOCK_DOMAIN_CROSSING;

  //====================================================================
  // Port Protocol Convertor / Data Width Convertor parameters
  //====================================================================
  parameter [1:0] MASTER0_TYPE  = 2'b10;      // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER1_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER2_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER3_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER4_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER5_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER6_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] MASTER7_TYPE  = MASTER0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3  
  
  parameter [1:0] SLAVE0_TYPE    = 2'b00;      // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE1_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE2_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE3_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE4_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE5_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE6_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE7_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3

  parameter [1:0] SLAVE8_TYPE      = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE9_TYPE      = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE10_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE11_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE12_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE13_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE14_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE15_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE16_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE17_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE18_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE19_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE20_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE21_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE22_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE23_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE24_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE25_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE26_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE27_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE28_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE29_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE30_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  parameter [1:0] SLAVE31_TYPE    = SLAVE0_TYPE;    // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3

  localparam [0:0] SLAVE0_READ_ZERO_SLAVE_ID    = 1'b1;                          // Disable slave read data interleave
  localparam [0:0] SLAVE1_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE2_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE3_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE4_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE5_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE6_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE7_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE8_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE9_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE10_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE11_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE12_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE13_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE14_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE15_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE16_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE17_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE18_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE19_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE20_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE21_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE22_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE23_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE24_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE25_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE26_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE27_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE28_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE29_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE30_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE31_READ_ZERO_SLAVE_ID    = SLAVE0_READ_ZERO_SLAVE_ID;    // Disable slave read data interleave

  localparam [0:0] SLAVE0_WRITE_ZERO_SLAVE_ID    = 1'b1;                           // Disable slave read data interleave
  localparam [0:0] SLAVE1_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE2_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE3_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE4_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE5_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE6_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE7_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;     // Disable slave read data interleave
  localparam [0:0] SLAVE8_WRITE_ZERO_SLAVE_ID     = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE9_WRITE_ZERO_SLAVE_ID     = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE10_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE11_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE12_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE13_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE14_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE15_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE16_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE17_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE18_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE19_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE20_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE21_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE22_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE23_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE24_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE25_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE26_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE27_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE28_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE29_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE30_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave
  localparam [0:0] SLAVE31_WRITE_ZERO_SLAVE_ID    = SLAVE0_WRITE_ZERO_SLAVE_ID;    // Disable slave read data interleave

  parameter  [1:0] AHB_MASTER0_BRESP_CHECK_MODE  =  2'b00;      // Defines wait response flag of Master0
  parameter  [1:0] AHB_MASTER1_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master1
  parameter  [1:0] AHB_MASTER2_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master2
  parameter  [1:0] AHB_MASTER3_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master3
  parameter  [1:0] AHB_MASTER4_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master4
  parameter  [1:0] AHB_MASTER5_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master5
  parameter  [1:0] AHB_MASTER6_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master6
  parameter  [1:0] AHB_MASTER7_BRESP_CHECK_MODE  =  AHB_MASTER0_BRESP_CHECK_MODE;      // Defines wait response flag of Master7
 
  parameter  [31:0] AHB_MASTER0_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER1_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER2_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER3_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER4_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER5_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER6_BRESP_CNT_WIDTH = 'h8;
  parameter  [31:0] AHB_MASTER7_BRESP_CNT_WIDTH = 'h8;

  parameter  [31:0] MASTER0_DATA_WIDTH  =  32;      // Defines data width of Master0
  parameter  [31:0] MASTER1_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master1
  parameter  [31:0] MASTER2_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master2
  parameter  [31:0] MASTER3_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master3
  parameter  [31:0] MASTER4_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master4
  parameter  [31:0] MASTER5_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master5
  parameter  [31:0] MASTER6_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master6
  parameter  [31:0] MASTER7_DATA_WIDTH  =  MASTER0_DATA_WIDTH;      // Defines data width of Master7
  
  parameter  [31:0] SLAVE0_DATA_WIDTH  =  32;      // Defines data width of Slave0
  parameter  [31:0] SLAVE1_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave1
  parameter  [31:0] SLAVE2_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave2
  parameter  [31:0] SLAVE3_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave3
  parameter  [31:0] SLAVE4_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave4
  parameter  [31:0] SLAVE5_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave5
  parameter  [31:0] SLAVE6_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave6
  parameter  [31:0] SLAVE7_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave7

  parameter  [31:0] SLAVE8_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave8
  parameter  [31:0] SLAVE9_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave9
  parameter  [31:0] SLAVE10_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave10
  parameter  [31:0] SLAVE11_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave11
  parameter  [31:0] SLAVE12_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave12
  parameter  [31:0] SLAVE13_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave13
  parameter  [31:0] SLAVE14_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave14
  parameter  [31:0] SLAVE15_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave15
  parameter  [31:0] SLAVE16_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave16
  parameter  [31:0] SLAVE17_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave17
  parameter  [31:0] SLAVE18_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave18
  parameter  [31:0] SLAVE19_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave19
  parameter  [31:0] SLAVE20_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave20
  parameter  [31:0] SLAVE21_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave21
  parameter  [31:0] SLAVE22_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave22
  parameter  [31:0] SLAVE23_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave23
  parameter  [31:0] SLAVE24_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave24
  parameter  [31:0] SLAVE25_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave25
  parameter  [31:0] SLAVE26_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave26
  parameter  [31:0] SLAVE27_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave27
  parameter  [31:0] SLAVE28_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave28
  parameter  [31:0] SLAVE29_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave29
  parameter  [31:0] SLAVE30_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave30
  parameter  [31:0] SLAVE31_DATA_WIDTH  =  SLAVE0_DATA_WIDTH;      // Defines data width of Slave31
  
  parameter integer  SLV_AXI4PRT_ADDRDEPTH = 2;          // Number transations width - 1 => 2 transations, 2 => 4 transations, etc.
  parameter integer  SLV_AXI4PRT_DATADEPTH = 2;          // Number transations width - 1 => 2 transations, 2 => 4 transations, etc.
  
  //====================================================================
  // Register Slice parameters
  //====================================================================
  parameter [0:0] MASTER0_CHAN_RS = 1'b1;
  parameter [0:0] MASTER1_CHAN_RS = MASTER0_CHAN_RS;
  parameter [0:0] MASTER2_CHAN_RS = MASTER0_CHAN_RS;
  parameter [0:0] MASTER3_CHAN_RS = MASTER0_CHAN_RS;
  parameter [0:0] MASTER4_CHAN_RS = MASTER0_CHAN_RS;
  parameter [0:0] MASTER5_CHAN_RS = MASTER0_CHAN_RS;
  parameter [0:0] MASTER6_CHAN_RS = MASTER0_CHAN_RS;
  parameter [0:0] MASTER7_CHAN_RS = MASTER0_CHAN_RS;
  
  parameter [0:0] SLAVE0_CHAN_RS = 1'b1;
  parameter [0:0] SLAVE1_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE2_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE3_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE4_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE5_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE6_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE7_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE8_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE9_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE10_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE11_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE12_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE13_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE14_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE15_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE16_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE17_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE18_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE19_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE20_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE21_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE22_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE23_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE24_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE25_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE26_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE27_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE28_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE29_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE30_CHAN_RS = SLAVE0_CHAN_RS;
  parameter [0:0] SLAVE31_CHAN_RS = SLAVE0_CHAN_RS;
  
  localparam [0:0]  MASTER0_AWCHAN_RS = MASTER0_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER1_AWCHAN_RS = MASTER1_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER2_AWCHAN_RS = MASTER2_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER3_AWCHAN_RS = MASTER3_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER4_AWCHAN_RS = MASTER4_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER5_AWCHAN_RS = MASTER5_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER6_AWCHAN_RS = MASTER6_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  MASTER7_AWCHAN_RS = MASTER7_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
              
  localparam [0:0]  MASTER0_ARCHAN_RS = MASTER0_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER1_ARCHAN_RS = MASTER1_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER2_ARCHAN_RS = MASTER2_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER3_ARCHAN_RS = MASTER3_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER4_ARCHAN_RS = MASTER4_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER5_ARCHAN_RS = MASTER5_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER6_ARCHAN_RS = MASTER6_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  MASTER7_ARCHAN_RS = MASTER7_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
             
  localparam [0:0]  MASTER0_WCHAN_RS = MASTER0_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER1_WCHAN_RS = MASTER1_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER2_WCHAN_RS = MASTER2_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER3_WCHAN_RS = MASTER3_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER4_WCHAN_RS = MASTER4_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER5_WCHAN_RS = MASTER5_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER6_WCHAN_RS = MASTER6_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  MASTER7_WCHAN_RS = MASTER7_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
             
  localparam [0:0]  MASTER0_RCHAN_RS = MASTER0_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER1_RCHAN_RS = MASTER1_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER2_RCHAN_RS = MASTER2_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER3_RCHAN_RS = MASTER3_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER4_RCHAN_RS = MASTER4_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER5_RCHAN_RS = MASTER5_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER6_RCHAN_RS = MASTER6_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  MASTER7_RCHAN_RS = MASTER7_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
              
  localparam [0:0]  MASTER0_BCHAN_RS = MASTER0_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER1_BCHAN_RS = MASTER1_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER2_BCHAN_RS = MASTER2_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER3_BCHAN_RS = MASTER3_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER4_BCHAN_RS = MASTER4_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER5_BCHAN_RS = MASTER5_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER6_BCHAN_RS = MASTER6_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  MASTER7_BCHAN_RS = MASTER7_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
              
  localparam [0:0]  SLAVE0_AWCHAN_RS  = SLAVE0_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE1_AWCHAN_RS  = SLAVE1_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE2_AWCHAN_RS  = SLAVE2_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE3_AWCHAN_RS  = SLAVE3_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE4_AWCHAN_RS  = SLAVE4_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE5_AWCHAN_RS  = SLAVE5_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE6_AWCHAN_RS  = SLAVE6_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE7_AWCHAN_RS  = SLAVE7_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE8_AWCHAN_RS  = SLAVE8_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE9_AWCHAN_RS  = SLAVE9_CHAN_RS;   // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE10_AWCHAN_RS = SLAVE10_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE11_AWCHAN_RS = SLAVE11_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE12_AWCHAN_RS = SLAVE12_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE13_AWCHAN_RS = SLAVE13_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE14_AWCHAN_RS = SLAVE14_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE15_AWCHAN_RS = SLAVE15_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE16_AWCHAN_RS = SLAVE16_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE17_AWCHAN_RS = SLAVE17_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE18_AWCHAN_RS = SLAVE18_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE19_AWCHAN_RS = SLAVE19_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE20_AWCHAN_RS = SLAVE20_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE21_AWCHAN_RS = SLAVE21_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE22_AWCHAN_RS = SLAVE22_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE23_AWCHAN_RS = SLAVE23_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE24_AWCHAN_RS = SLAVE24_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE25_AWCHAN_RS = SLAVE25_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE26_AWCHAN_RS = SLAVE26_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE27_AWCHAN_RS = SLAVE27_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE28_AWCHAN_RS = SLAVE28_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE29_AWCHAN_RS = SLAVE29_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE30_AWCHAN_RS = SLAVE30_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [0:0]  SLAVE31_AWCHAN_RS = SLAVE31_CHAN_RS;  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
              
  localparam [0:0]  SLAVE0_ARCHAN_RS  = SLAVE0_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE1_ARCHAN_RS  = SLAVE1_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE2_ARCHAN_RS  = SLAVE2_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE3_ARCHAN_RS  = SLAVE3_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE4_ARCHAN_RS  = SLAVE4_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE5_ARCHAN_RS  = SLAVE5_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE6_ARCHAN_RS  = SLAVE6_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE7_ARCHAN_RS  = SLAVE7_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE8_ARCHAN_RS  = SLAVE8_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE9_ARCHAN_RS  = SLAVE9_CHAN_RS;   // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE10_ARCHAN_RS = SLAVE10_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE11_ARCHAN_RS = SLAVE11_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE12_ARCHAN_RS = SLAVE12_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE13_ARCHAN_RS = SLAVE13_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE14_ARCHAN_RS = SLAVE14_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE15_ARCHAN_RS = SLAVE15_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE16_ARCHAN_RS = SLAVE16_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE17_ARCHAN_RS = SLAVE17_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE18_ARCHAN_RS = SLAVE18_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE19_ARCHAN_RS = SLAVE19_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE20_ARCHAN_RS = SLAVE20_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE21_ARCHAN_RS = SLAVE21_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE22_ARCHAN_RS = SLAVE22_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE23_ARCHAN_RS = SLAVE23_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE24_ARCHAN_RS = SLAVE24_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE25_ARCHAN_RS = SLAVE25_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE26_ARCHAN_RS = SLAVE26_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE27_ARCHAN_RS = SLAVE27_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE28_ARCHAN_RS = SLAVE28_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE29_ARCHAN_RS = SLAVE29_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE30_ARCHAN_RS = SLAVE30_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [0:0]  SLAVE31_ARCHAN_RS = SLAVE31_CHAN_RS;  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  
  localparam [0:0]  SLAVE0_WCHAN_RS  = SLAVE0_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE1_WCHAN_RS  = SLAVE1_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE2_WCHAN_RS  = SLAVE2_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE3_WCHAN_RS  = SLAVE3_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE4_WCHAN_RS  = SLAVE4_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE5_WCHAN_RS  = SLAVE5_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE6_WCHAN_RS  = SLAVE6_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE7_WCHAN_RS  = SLAVE7_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE8_WCHAN_RS  = SLAVE8_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE9_WCHAN_RS  = SLAVE9_CHAN_RS;   // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE10_WCHAN_RS = SLAVE10_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE11_WCHAN_RS = SLAVE11_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE12_WCHAN_RS = SLAVE12_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE13_WCHAN_RS = SLAVE13_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE14_WCHAN_RS = SLAVE14_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE15_WCHAN_RS = SLAVE15_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE16_WCHAN_RS = SLAVE16_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE17_WCHAN_RS = SLAVE17_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE18_WCHAN_RS = SLAVE18_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE19_WCHAN_RS = SLAVE19_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE20_WCHAN_RS = SLAVE20_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE21_WCHAN_RS = SLAVE21_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE22_WCHAN_RS = SLAVE22_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE23_WCHAN_RS = SLAVE23_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE24_WCHAN_RS = SLAVE24_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE25_WCHAN_RS = SLAVE25_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE26_WCHAN_RS = SLAVE26_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE27_WCHAN_RS = SLAVE27_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE28_WCHAN_RS = SLAVE28_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE29_WCHAN_RS = SLAVE29_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE30_WCHAN_RS = SLAVE30_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [0:0]  SLAVE31_WCHAN_RS = SLAVE31_CHAN_RS;  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  
  localparam [0:0]  SLAVE0_RCHAN_RS  = SLAVE0_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE1_RCHAN_RS  = SLAVE1_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE2_RCHAN_RS  = SLAVE2_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE3_RCHAN_RS  = SLAVE3_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE4_RCHAN_RS  = SLAVE4_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE5_RCHAN_RS  = SLAVE5_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE6_RCHAN_RS  = SLAVE6_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE7_RCHAN_RS  = SLAVE7_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE8_RCHAN_RS  = SLAVE8_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE9_RCHAN_RS  = SLAVE9_CHAN_RS;   // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE10_RCHAN_RS = SLAVE10_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE11_RCHAN_RS = SLAVE11_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE12_RCHAN_RS = SLAVE12_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE13_RCHAN_RS = SLAVE13_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE14_RCHAN_RS = SLAVE14_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE15_RCHAN_RS = SLAVE15_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE16_RCHAN_RS = SLAVE16_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE17_RCHAN_RS = SLAVE17_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE18_RCHAN_RS = SLAVE18_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE19_RCHAN_RS = SLAVE19_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE20_RCHAN_RS = SLAVE20_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE21_RCHAN_RS = SLAVE21_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE22_RCHAN_RS = SLAVE22_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE23_RCHAN_RS = SLAVE23_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE24_RCHAN_RS = SLAVE24_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE25_RCHAN_RS = SLAVE25_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE26_RCHAN_RS = SLAVE26_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE27_RCHAN_RS = SLAVE27_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE28_RCHAN_RS = SLAVE28_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE29_RCHAN_RS = SLAVE29_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE30_RCHAN_RS = SLAVE30_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [0:0]  SLAVE31_RCHAN_RS = SLAVE31_CHAN_RS;  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  
  localparam [0:0]  SLAVE0_BCHAN_RS  = SLAVE0_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE1_BCHAN_RS  = SLAVE1_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE2_BCHAN_RS  = SLAVE2_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE3_BCHAN_RS  = SLAVE3_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE4_BCHAN_RS  = SLAVE4_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE5_BCHAN_RS  = SLAVE5_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE6_BCHAN_RS  = SLAVE6_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE7_BCHAN_RS  = SLAVE7_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE8_BCHAN_RS  = SLAVE8_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE9_BCHAN_RS  = SLAVE9_CHAN_RS;   // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE10_BCHAN_RS = SLAVE10_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE11_BCHAN_RS = SLAVE11_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE12_BCHAN_RS = SLAVE12_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE13_BCHAN_RS = SLAVE13_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE14_BCHAN_RS = SLAVE14_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE15_BCHAN_RS = SLAVE15_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE16_BCHAN_RS = SLAVE16_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE17_BCHAN_RS = SLAVE17_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE18_BCHAN_RS = SLAVE18_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE19_BCHAN_RS = SLAVE19_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE20_BCHAN_RS = SLAVE20_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE21_BCHAN_RS = SLAVE21_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE22_BCHAN_RS = SLAVE22_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE23_BCHAN_RS = SLAVE23_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE24_BCHAN_RS = SLAVE24_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE25_BCHAN_RS = SLAVE25_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE26_BCHAN_RS = SLAVE26_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE27_BCHAN_RS = SLAVE27_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE28_BCHAN_RS = SLAVE28_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE29_BCHAN_RS = SLAVE29_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE30_BCHAN_RS = SLAVE30_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [0:0]  SLAVE31_BCHAN_RS = SLAVE31_CHAN_RS;  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  
     //===================================================================================================================================


  parameter  [7:0] MASTER0_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master0
  parameter  [7:0] MASTER1_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master1
  parameter  [7:0] MASTER2_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master2
  parameter  [7:0] MASTER3_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master3
  parameter  [7:0] MASTER4_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master4
  parameter  [7:0] MASTER5_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master5
  parameter  [7:0] MASTER6_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master6
  parameter  [7:0] MASTER7_DEF_BURST_LEN  =  8'h0;      // Defines the default burst length if the AHB interface of Master7

  parameter  [13:0] SLAVE0_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave0
  parameter  [13:0] SLAVE1_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave1
  parameter  [13:0] SLAVE2_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave2
  parameter  [13:0] SLAVE3_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave3
  parameter  [13:0] SLAVE4_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave4
  parameter  [13:0] SLAVE5_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave5
  parameter  [13:0] SLAVE6_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave6
  parameter  [13:0] SLAVE7_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave7
  
  parameter  [13:0] SLAVE8_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave8
  parameter  [13:0] SLAVE9_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave9
  parameter  [13:0] SLAVE10_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave10
  parameter  [13:0] SLAVE11_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave11
  parameter  [13:0] SLAVE12_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave12
  parameter  [13:0] SLAVE13_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave13
  parameter  [13:0] SLAVE14_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave14
  parameter  [13:0] SLAVE15_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave15
  parameter  [13:0] SLAVE16_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave16
  parameter  [13:0] SLAVE17_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave17
  parameter  [13:0] SLAVE18_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave18
  parameter  [13:0] SLAVE19_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave19
  parameter  [13:0] SLAVE20_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave20
  parameter  [13:0] SLAVE21_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave21
  parameter  [13:0] SLAVE22_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave22
  parameter  [13:0] SLAVE23_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave23
  parameter  [13:0] SLAVE24_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave24
  parameter  [13:0] SLAVE25_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave25
  parameter  [13:0] SLAVE26_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave26
  parameter  [13:0] SLAVE27_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave27
  parameter  [13:0] SLAVE28_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave28
  parameter  [13:0] SLAVE29_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave29
  parameter  [13:0] SLAVE30_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave30
  parameter  [13:0] SLAVE31_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Slave31

  
  parameter  [13:0] MASTER0_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master0
  parameter  [13:0] MASTER1_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master1
  parameter  [13:0] MASTER2_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master2
  parameter  [13:0] MASTER3_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master3
  parameter  [13:0] MASTER4_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master4
  parameter  [13:0] MASTER5_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master5
  parameter  [13:0] MASTER6_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master6
  parameter  [13:0] MASTER7_DWC_DATA_FIFO_DEPTH  =  14'h10;      // Defines the depth of the data caxi4interconnect_FIFO in the datawidth converter of Master7

  parameter integer DWC_ADDR_FIFO_DEPTH_CEILING = 'h10;

  parameter integer NUM_MASTERS_WIDTH  = (NUM_MASTERS == 1) ? 1 : $clog2(NUM_MASTERS);
  
  localparam HI_FREQ = ((CROSSBAR_MODE == 1) || ((CROSSBAR_MODE == 0) && (RD_ARB_EN == 0))) ? 1 : 0;        // increases freq of operation at cost of added latency
  
  localparam integer NUM_SLAVES_WIDTH  = (NUM_SLAVES == 1) ? 1 : $clog2(NUM_SLAVES);
            
  localparam integer ADDR_WIDTH_BITS  = ( ADDR_WIDTH <= 16 ) ? 4 : $clog2(ADDR_WIDTH);

  localparam NUM_THREADS_WIDTH    =  (NUM_THREADS == 1) ? 1 : $clog2(NUM_THREADS);

  localparam OPEN_TRANS_WIDTH    = ( OPEN_TRANS_MAX == 1 ) ? 1 : $clog2(OPEN_TRANS_MAX);
    
  localparam MASTERID_WIDTH    = ( NUM_MASTERS_WIDTH + ID_WIDTH );      // defines width masterID - includes infrastructure port number plus ID
  
  localparam  BASE_WIDTH = ADDR_WIDTH;//-UPPER_COMPARE_BIT;

  localparam [ ( NUM_SLAVES* BASE_WIDTH )-1 : 0 ]   SLOT_BASE_VEC = { SLOT31_BASE_VEC[BASE_WIDTH-1:0], SLOT30_BASE_VEC[BASE_WIDTH-1:0], SLOT29_BASE_VEC[BASE_WIDTH-1:0], SLOT28_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT27_BASE_VEC[BASE_WIDTH-1:0], SLOT26_BASE_VEC[BASE_WIDTH-1:0], SLOT25_BASE_VEC[BASE_WIDTH-1:0], SLOT24_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT23_BASE_VEC[BASE_WIDTH-1:0], SLOT22_BASE_VEC[BASE_WIDTH-1:0], SLOT21_BASE_VEC[BASE_WIDTH-1:0], SLOT20_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT19_BASE_VEC[BASE_WIDTH-1:0], SLOT18_BASE_VEC[BASE_WIDTH-1:0], SLOT17_BASE_VEC[BASE_WIDTH-1:0], SLOT16_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT15_BASE_VEC[BASE_WIDTH-1:0], SLOT14_BASE_VEC[BASE_WIDTH-1:0], SLOT13_BASE_VEC[BASE_WIDTH-1:0], SLOT12_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT11_BASE_VEC[BASE_WIDTH-1:0], SLOT10_BASE_VEC[BASE_WIDTH-1:0], SLOT9_BASE_VEC[BASE_WIDTH-1:0], SLOT8_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT7_BASE_VEC[BASE_WIDTH-1:0], SLOT6_BASE_VEC[BASE_WIDTH-1:0], SLOT5_BASE_VEC[BASE_WIDTH-1:0], SLOT4_BASE_VEC[BASE_WIDTH-1:0],
                                                                      SLOT3_BASE_VEC[BASE_WIDTH-1:0], SLOT2_BASE_VEC[BASE_WIDTH-1:0], SLOT1_BASE_VEC[BASE_WIDTH-1:0], SLOT0_BASE_VEC[BASE_WIDTH-1:0] };
                                                          

  
  localparam CMPR_WIDTH = UPPER_COMPARE_BIT-LOWER_COMPARE_BIT;

  localparam [ ( NUM_SLAVES* (CMPR_WIDTH) )-1 : 0 ]   SLOT_MIN_VEC  = 
                              { SLOT31_MIN_VEC[CMPR_WIDTH-1:0], SLOT30_MIN_VEC[CMPR_WIDTH-1:0], SLOT29_MIN_VEC[CMPR_WIDTH-1:0], SLOT28_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT27_MIN_VEC[CMPR_WIDTH-1:0], SLOT26_MIN_VEC[CMPR_WIDTH-1:0], SLOT25_MIN_VEC[CMPR_WIDTH-1:0], SLOT24_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT23_MIN_VEC[CMPR_WIDTH-1:0], SLOT22_MIN_VEC[CMPR_WIDTH-1:0], SLOT21_MIN_VEC[CMPR_WIDTH-1:0], SLOT20_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT19_MIN_VEC[CMPR_WIDTH-1:0], SLOT18_MIN_VEC[CMPR_WIDTH-1:0], SLOT17_MIN_VEC[CMPR_WIDTH-1:0], SLOT16_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT15_MIN_VEC[CMPR_WIDTH-1:0], SLOT14_MIN_VEC[CMPR_WIDTH-1:0], SLOT13_MIN_VEC[CMPR_WIDTH-1:0], SLOT12_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT11_MIN_VEC[CMPR_WIDTH-1:0], SLOT10_MIN_VEC[CMPR_WIDTH-1:0], SLOT9_MIN_VEC[CMPR_WIDTH-1:0],  SLOT8_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT7_MIN_VEC[CMPR_WIDTH-1:0],  SLOT6_MIN_VEC[CMPR_WIDTH-1:0],  SLOT5_MIN_VEC[CMPR_WIDTH-1:0],  SLOT4_MIN_VEC[CMPR_WIDTH-1:0],
                                SLOT3_MIN_VEC[CMPR_WIDTH-1:0],  SLOT2_MIN_VEC[CMPR_WIDTH-1:0],  SLOT1_MIN_VEC[CMPR_WIDTH-1:0],  SLOT0_MIN_VEC[CMPR_WIDTH-1:0] };        // SLOT Min per slave 
                            
  localparam [ ( NUM_SLAVES* (CMPR_WIDTH) )-1 : 0 ]   SLOT_MAX_VEC  = 
                              { SLOT31_MAX_VEC[CMPR_WIDTH-1:0], SLOT30_MAX_VEC[CMPR_WIDTH-1:0], SLOT29_MAX_VEC[CMPR_WIDTH-1:0], SLOT28_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT27_MAX_VEC[CMPR_WIDTH-1:0], SLOT26_MAX_VEC[CMPR_WIDTH-1:0], SLOT25_MAX_VEC[CMPR_WIDTH-1:0], SLOT24_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT23_MAX_VEC[CMPR_WIDTH-1:0], SLOT22_MAX_VEC[CMPR_WIDTH-1:0], SLOT21_MAX_VEC[CMPR_WIDTH-1:0], SLOT20_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT19_MAX_VEC[CMPR_WIDTH-1:0], SLOT18_MAX_VEC[CMPR_WIDTH-1:0], SLOT17_MAX_VEC[CMPR_WIDTH-1:0], SLOT16_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT15_MAX_VEC[CMPR_WIDTH-1:0], SLOT14_MAX_VEC[CMPR_WIDTH-1:0], SLOT13_MAX_VEC[CMPR_WIDTH-1:0], SLOT12_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT11_MAX_VEC[CMPR_WIDTH-1:0], SLOT10_MAX_VEC[CMPR_WIDTH-1:0], SLOT9_MAX_VEC[CMPR_WIDTH-1:0],  SLOT8_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT7_MAX_VEC[CMPR_WIDTH-1:0],  SLOT6_MAX_VEC[CMPR_WIDTH-1:0],  SLOT5_MAX_VEC[CMPR_WIDTH-1:0],  SLOT4_MAX_VEC[CMPR_WIDTH-1:0],
                                SLOT3_MAX_VEC[CMPR_WIDTH-1:0],  SLOT2_MAX_VEC[CMPR_WIDTH-1:0],  SLOT1_MAX_VEC[CMPR_WIDTH-1:0],  SLOT0_MAX_VEC[CMPR_WIDTH-1:0] };        // SLOT Max per slave
                                
  // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3, 10 = AHB
  localparam [(NUM_MASTERS*2)-1:0] MASTER_TYPE  = { MASTER7_TYPE, MASTER6_TYPE, MASTER5_TYPE, MASTER4_TYPE,
                                                    MASTER3_TYPE, MASTER2_TYPE, MASTER1_TYPE, MASTER0_TYPE };    
  
  //SAR76987 SMG should be NUM_SLAVES not NUM_MASTERS
  // Valid Values - 00 = AXI4, 01=AXI4-Lite, 11 = AXI3
  localparam [(NUM_SLAVES*2)-1:0] SLAVE_TYPE    = { SLAVE31_TYPE, SLAVE30_TYPE, SLAVE29_TYPE, SLAVE28_TYPE, SLAVE27_TYPE, SLAVE26_TYPE, SLAVE25_TYPE, SLAVE24_TYPE,
                                                    SLAVE23_TYPE, SLAVE22_TYPE, SLAVE21_TYPE, SLAVE20_TYPE, SLAVE19_TYPE, SLAVE18_TYPE, SLAVE17_TYPE, SLAVE16_TYPE,
                                                    SLAVE15_TYPE, SLAVE14_TYPE, SLAVE13_TYPE, SLAVE12_TYPE, SLAVE11_TYPE, SLAVE10_TYPE, SLAVE9_TYPE,  SLAVE8_TYPE,
                                                    SLAVE7_TYPE,  SLAVE6_TYPE,  SLAVE5_TYPE,  SLAVE4_TYPE,  SLAVE3_TYPE,  SLAVE2_TYPE,  SLAVE1_TYPE,  SLAVE0_TYPE };    

  localparam [NUM_SLAVES-1:0] SLAVE_READ_ZERO_SLAVE_ID    = { SLAVE31_READ_ZERO_SLAVE_ID, SLAVE30_READ_ZERO_SLAVE_ID, SLAVE29_READ_ZERO_SLAVE_ID, SLAVE28_READ_ZERO_SLAVE_ID, SLAVE27_READ_ZERO_SLAVE_ID, SLAVE26_READ_ZERO_SLAVE_ID, SLAVE25_READ_ZERO_SLAVE_ID, SLAVE24_READ_ZERO_SLAVE_ID,
                                                    SLAVE23_READ_ZERO_SLAVE_ID, SLAVE22_READ_ZERO_SLAVE_ID, SLAVE21_READ_ZERO_SLAVE_ID, SLAVE20_READ_ZERO_SLAVE_ID, SLAVE19_READ_ZERO_SLAVE_ID, SLAVE18_READ_ZERO_SLAVE_ID, SLAVE17_READ_ZERO_SLAVE_ID, SLAVE16_READ_ZERO_SLAVE_ID,
                                                    SLAVE15_READ_ZERO_SLAVE_ID, SLAVE14_READ_ZERO_SLAVE_ID, SLAVE13_READ_ZERO_SLAVE_ID, SLAVE12_READ_ZERO_SLAVE_ID, SLAVE11_READ_ZERO_SLAVE_ID, SLAVE10_READ_ZERO_SLAVE_ID, SLAVE9_READ_ZERO_SLAVE_ID,  SLAVE8_READ_ZERO_SLAVE_ID,
                                                    SLAVE7_READ_ZERO_SLAVE_ID,  SLAVE6_READ_ZERO_SLAVE_ID,  SLAVE5_READ_ZERO_SLAVE_ID,  SLAVE4_READ_ZERO_SLAVE_ID,  SLAVE3_READ_ZERO_SLAVE_ID,  SLAVE2_READ_ZERO_SLAVE_ID,  SLAVE1_READ_ZERO_SLAVE_ID,  SLAVE0_READ_ZERO_SLAVE_ID };    

  localparam [NUM_SLAVES-1:0] SLAVE_WRITE_ZERO_SLAVE_ID    = { SLAVE31_WRITE_ZERO_SLAVE_ID, SLAVE30_WRITE_ZERO_SLAVE_ID, SLAVE29_WRITE_ZERO_SLAVE_ID, SLAVE28_WRITE_ZERO_SLAVE_ID, SLAVE27_WRITE_ZERO_SLAVE_ID, SLAVE26_WRITE_ZERO_SLAVE_ID, SLAVE25_WRITE_ZERO_SLAVE_ID, SLAVE24_WRITE_ZERO_SLAVE_ID,
                                                    SLAVE23_WRITE_ZERO_SLAVE_ID, SLAVE22_WRITE_ZERO_SLAVE_ID, SLAVE21_WRITE_ZERO_SLAVE_ID, SLAVE20_WRITE_ZERO_SLAVE_ID, SLAVE19_WRITE_ZERO_SLAVE_ID, SLAVE18_WRITE_ZERO_SLAVE_ID, SLAVE17_WRITE_ZERO_SLAVE_ID, SLAVE16_WRITE_ZERO_SLAVE_ID,
                                                    SLAVE15_WRITE_ZERO_SLAVE_ID, SLAVE14_WRITE_ZERO_SLAVE_ID, SLAVE13_WRITE_ZERO_SLAVE_ID, SLAVE12_WRITE_ZERO_SLAVE_ID, SLAVE11_WRITE_ZERO_SLAVE_ID, SLAVE10_WRITE_ZERO_SLAVE_ID, SLAVE9_WRITE_ZERO_SLAVE_ID,  SLAVE8_WRITE_ZERO_SLAVE_ID,
                                                    SLAVE7_WRITE_ZERO_SLAVE_ID,  SLAVE6_WRITE_ZERO_SLAVE_ID,  SLAVE5_WRITE_ZERO_SLAVE_ID,  SLAVE4_WRITE_ZERO_SLAVE_ID,  SLAVE3_WRITE_ZERO_SLAVE_ID,  SLAVE2_WRITE_ZERO_SLAVE_ID,  SLAVE1_WRITE_ZERO_SLAVE_ID,  SLAVE0_WRITE_ZERO_SLAVE_ID };    

  localparam [NUM_MASTERS-1:0]  MASTER_AWCHAN_RS = { MASTER7_AWCHAN_RS, MASTER6_AWCHAN_RS, MASTER5_AWCHAN_RS, MASTER4_AWCHAN_RS,  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
                                                    MASTER3_AWCHAN_RS, MASTER2_AWCHAN_RS, MASTER1_AWCHAN_RS, MASTER0_AWCHAN_RS };

  localparam [NUM_MASTERS-1:0]  MASTER_ARCHAN_RS = { MASTER7_ARCHAN_RS, MASTER6_ARCHAN_RS, MASTER5_ARCHAN_RS, MASTER4_ARCHAN_RS,  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
                                                    MASTER3_ARCHAN_RS, MASTER2_ARCHAN_RS, MASTER1_ARCHAN_RS, MASTER0_ARCHAN_RS };

  localparam [NUM_MASTERS-1:0]  MASTER_WCHAN_RS = { MASTER7_WCHAN_RS, MASTER6_WCHAN_RS, MASTER5_WCHAN_RS, MASTER4_WCHAN_RS,    // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
                                                    MASTER3_WCHAN_RS, MASTER2_WCHAN_RS, MASTER1_WCHAN_RS, MASTER0_WCHAN_RS };

  localparam [NUM_MASTERS-1:0]  MASTER_RCHAN_RS = { MASTER7_RCHAN_RS, MASTER6_RCHAN_RS, MASTER5_RCHAN_RS, MASTER4_RCHAN_RS,    // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
                                                    MASTER3_RCHAN_RS, MASTER2_RCHAN_RS, MASTER1_RCHAN_RS, MASTER0_RCHAN_RS };

  localparam [NUM_MASTERS-1:0]  MASTER_BCHAN_RS = { MASTER7_BCHAN_RS, MASTER6_BCHAN_RS, MASTER5_BCHAN_RS, MASTER4_BCHAN_RS,    // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
                                                    MASTER3_BCHAN_RS, MASTER2_BCHAN_RS, MASTER1_BCHAN_RS, MASTER0_BCHAN_RS };

                                                    
  // 0 - no AWCHAN register slice, 1 - AWCHAN register slice inserted
  localparam [NUM_SLAVES-1:0] SLAVE_AWCHAN_RS = { SLAVE31_AWCHAN_RS, SLAVE30_AWCHAN_RS, SLAVE29_AWCHAN_RS, SLAVE28_AWCHAN_RS, SLAVE27_AWCHAN_RS, SLAVE26_AWCHAN_RS, SLAVE25_AWCHAN_RS, SLAVE24_AWCHAN_RS,
                                                  SLAVE23_AWCHAN_RS, SLAVE22_AWCHAN_RS, SLAVE21_AWCHAN_RS, SLAVE20_AWCHAN_RS, SLAVE19_AWCHAN_RS, SLAVE18_AWCHAN_RS, SLAVE17_AWCHAN_RS, SLAVE16_AWCHAN_RS,
                                                  SLAVE15_AWCHAN_RS, SLAVE14_AWCHAN_RS, SLAVE13_AWCHAN_RS, SLAVE12_AWCHAN_RS, SLAVE11_AWCHAN_RS, SLAVE10_AWCHAN_RS, SLAVE9_AWCHAN_RS,  SLAVE8_AWCHAN_RS,
                                                  SLAVE7_AWCHAN_RS,  SLAVE6_AWCHAN_RS,  SLAVE5_AWCHAN_RS,  SLAVE4_AWCHAN_RS,  SLAVE3_AWCHAN_RS,  SLAVE2_AWCHAN_RS,  SLAVE1_AWCHAN_RS,  SLAVE0_AWCHAN_RS };
  
  // 0 - no ARCHAN register slice, 1 - ARCHAN register slice inserted
  localparam [NUM_SLAVES-1:0] SLAVE_ARCHAN_RS = { SLAVE31_ARCHAN_RS, SLAVE30_ARCHAN_RS, SLAVE29_ARCHAN_RS, SLAVE28_ARCHAN_RS, SLAVE27_ARCHAN_RS, SLAVE26_ARCHAN_RS, SLAVE25_ARCHAN_RS, SLAVE24_ARCHAN_RS,
                                                  SLAVE23_ARCHAN_RS, SLAVE22_ARCHAN_RS, SLAVE21_ARCHAN_RS, SLAVE20_ARCHAN_RS, SLAVE19_ARCHAN_RS, SLAVE18_ARCHAN_RS, SLAVE17_ARCHAN_RS, SLAVE16_ARCHAN_RS,
                                                  SLAVE15_ARCHAN_RS, SLAVE14_ARCHAN_RS, SLAVE13_ARCHAN_RS, SLAVE12_ARCHAN_RS, SLAVE11_ARCHAN_RS, SLAVE10_ARCHAN_RS, SLAVE9_ARCHAN_RS,  SLAVE8_ARCHAN_RS,
                                                  SLAVE7_ARCHAN_RS,  SLAVE6_ARCHAN_RS,  SLAVE5_ARCHAN_RS,  SLAVE4_ARCHAN_RS,  SLAVE3_ARCHAN_RS,  SLAVE2_ARCHAN_RS,  SLAVE1_ARCHAN_RS,  SLAVE0_ARCHAN_RS };

  // 0 - no WCHAN register slice, 1 - WCHAN register slice inserted
  localparam [NUM_SLAVES-1:0] SLAVE_WCHAN_RS = { SLAVE31_WCHAN_RS, SLAVE30_WCHAN_RS, SLAVE29_WCHAN_RS, SLAVE28_WCHAN_RS, SLAVE27_WCHAN_RS, SLAVE26_WCHAN_RS, SLAVE25_WCHAN_RS, SLAVE24_WCHAN_RS,
                                                 SLAVE23_WCHAN_RS, SLAVE22_WCHAN_RS, SLAVE21_WCHAN_RS, SLAVE20_WCHAN_RS, SLAVE19_WCHAN_RS, SLAVE18_WCHAN_RS, SLAVE17_WCHAN_RS, SLAVE16_WCHAN_RS,
                                                 SLAVE15_WCHAN_RS, SLAVE14_WCHAN_RS, SLAVE13_WCHAN_RS, SLAVE12_WCHAN_RS, SLAVE11_WCHAN_RS, SLAVE10_WCHAN_RS, SLAVE9_WCHAN_RS,  SLAVE8_WCHAN_RS,
                                                 SLAVE7_WCHAN_RS,  SLAVE6_WCHAN_RS,  SLAVE5_WCHAN_RS,  SLAVE4_WCHAN_RS,  SLAVE3_WCHAN_RS,  SLAVE2_WCHAN_RS,  SLAVE1_WCHAN_RS,  SLAVE0_WCHAN_RS  };

  // 0 - no RCHAN register slice, 1 - RCHAN register slice inserted
  localparam [NUM_SLAVES-1:0] SLAVE_RCHAN_RS = { SLAVE31_RCHAN_RS, SLAVE30_RCHAN_RS, SLAVE29_RCHAN_RS, SLAVE28_RCHAN_RS, SLAVE27_RCHAN_RS, SLAVE26_RCHAN_RS, SLAVE25_RCHAN_RS, SLAVE24_RCHAN_RS,
                                                 SLAVE23_RCHAN_RS, SLAVE22_RCHAN_RS, SLAVE21_RCHAN_RS, SLAVE20_RCHAN_RS, SLAVE19_RCHAN_RS, SLAVE18_RCHAN_RS, SLAVE17_RCHAN_RS, SLAVE16_RCHAN_RS,
                                                 SLAVE15_RCHAN_RS, SLAVE14_RCHAN_RS, SLAVE13_RCHAN_RS, SLAVE12_RCHAN_RS, SLAVE11_RCHAN_RS, SLAVE10_RCHAN_RS, SLAVE9_RCHAN_RS,  SLAVE8_RCHAN_RS,
                                                 SLAVE7_RCHAN_RS,  SLAVE6_RCHAN_RS,  SLAVE5_RCHAN_RS,  SLAVE4_RCHAN_RS,  SLAVE3_RCHAN_RS,  SLAVE2_RCHAN_RS,  SLAVE1_RCHAN_RS,  SLAVE0_RCHAN_RS  };

  // 0 - no BCHAN register slice, 1 - BCHAN register slice inserted
  localparam [NUM_SLAVES-1:0] SLAVE_BCHAN_RS = { SLAVE31_BCHAN_RS, SLAVE30_BCHAN_RS, SLAVE29_BCHAN_RS, SLAVE28_BCHAN_RS, SLAVE27_BCHAN_RS, SLAVE26_BCHAN_RS, SLAVE25_BCHAN_RS, SLAVE24_BCHAN_RS,
                                                 SLAVE23_BCHAN_RS, SLAVE22_BCHAN_RS, SLAVE21_BCHAN_RS, SLAVE20_BCHAN_RS, SLAVE19_BCHAN_RS, SLAVE18_BCHAN_RS, SLAVE17_BCHAN_RS, SLAVE16_BCHAN_RS,
                                                 SLAVE15_BCHAN_RS, SLAVE14_BCHAN_RS, SLAVE13_BCHAN_RS, SLAVE12_BCHAN_RS, SLAVE11_BCHAN_RS, SLAVE10_BCHAN_RS, SLAVE9_BCHAN_RS,  SLAVE8_BCHAN_RS,
                                                 SLAVE7_BCHAN_RS,  SLAVE6_BCHAN_RS,  SLAVE5_BCHAN_RS,  SLAVE4_BCHAN_RS,  SLAVE3_BCHAN_RS,  SLAVE2_BCHAN_RS,  SLAVE1_BCHAN_RS,  SLAVE0_BCHAN_RS };

  localparam [(2*NUM_MASTERS)-1:0] AHB_MASTER_PORTS_BRESP_CHECK_MODE = { AHB_MASTER7_BRESP_CHECK_MODE,
                                      AHB_MASTER6_BRESP_CHECK_MODE,
                                      AHB_MASTER5_BRESP_CHECK_MODE,
                                      AHB_MASTER4_BRESP_CHECK_MODE,
                                      AHB_MASTER3_BRESP_CHECK_MODE,
                                      AHB_MASTER2_BRESP_CHECK_MODE,
                                      AHB_MASTER1_BRESP_CHECK_MODE,
                                      AHB_MASTER0_BRESP_CHECK_MODE
                                      };

  localparam [(32*NUM_MASTERS)-1:0] AHB_MASTER_PORTS_BRESP_CNT_WIDTH = { AHB_MASTER7_BRESP_CNT_WIDTH,
                                      AHB_MASTER6_BRESP_CNT_WIDTH,
                                      AHB_MASTER5_BRESP_CNT_WIDTH,
                                      AHB_MASTER4_BRESP_CNT_WIDTH,
                                      AHB_MASTER3_BRESP_CNT_WIDTH,
                                      AHB_MASTER2_BRESP_CNT_WIDTH,
                                      AHB_MASTER1_BRESP_CNT_WIDTH,
                                      AHB_MASTER0_BRESP_CNT_WIDTH
                                      };



  localparam [(NUM_MASTERS*32)-1:0] MASTER_PORTS_DATA_WIDTH = { MASTER7_DATA_WIDTH,
                                      MASTER6_DATA_WIDTH,
                                      MASTER5_DATA_WIDTH,
                                      MASTER4_DATA_WIDTH,
                                      MASTER3_DATA_WIDTH,
                                      MASTER2_DATA_WIDTH,
                                      MASTER1_DATA_WIDTH,
                                      MASTER0_DATA_WIDTH
                                      };
  
  localparam [(NUM_SLAVES*32)-1:0]  SLAVE_PORTS_DATA_WIDTH  = 
                                      {
                                      SLAVE31_DATA_WIDTH,
                                      SLAVE30_DATA_WIDTH,
                                      SLAVE29_DATA_WIDTH,
                                      SLAVE28_DATA_WIDTH,
                                      SLAVE27_DATA_WIDTH,
                                      SLAVE26_DATA_WIDTH,
                                      SLAVE25_DATA_WIDTH,
                                      SLAVE24_DATA_WIDTH,
                                      SLAVE23_DATA_WIDTH,
                                      SLAVE22_DATA_WIDTH,
                                      SLAVE21_DATA_WIDTH,
                                      SLAVE20_DATA_WIDTH,
                                      SLAVE19_DATA_WIDTH,
                                      SLAVE18_DATA_WIDTH,
                                      SLAVE17_DATA_WIDTH,
                                      SLAVE16_DATA_WIDTH,  
                                      SLAVE15_DATA_WIDTH,
                                      SLAVE14_DATA_WIDTH,
                                      SLAVE13_DATA_WIDTH,
                                      SLAVE12_DATA_WIDTH,
                                      SLAVE11_DATA_WIDTH,
                                      SLAVE10_DATA_WIDTH,
                                      SLAVE9_DATA_WIDTH,
                                      SLAVE8_DATA_WIDTH,
                                      SLAVE7_DATA_WIDTH,
                                      SLAVE6_DATA_WIDTH,
                                      SLAVE5_DATA_WIDTH,
                                      SLAVE4_DATA_WIDTH,
                                      SLAVE3_DATA_WIDTH,
                                      SLAVE2_DATA_WIDTH,
                                      SLAVE1_DATA_WIDTH,
                                      SLAVE0_DATA_WIDTH
                                      };
                          
                                    
  localparam integer MASTER_DATA_WIDTH_PORT = ( MASTER7_DATA_WIDTH + MASTER6_DATA_WIDTH + MASTER5_DATA_WIDTH + MASTER4_DATA_WIDTH + 
                                                MASTER3_DATA_WIDTH + MASTER2_DATA_WIDTH + MASTER1_DATA_WIDTH + MASTER0_DATA_WIDTH);
  
  localparam [12:0] MDW0_UPPER = MASTER0_DATA_WIDTH;
  localparam [12:0] MDW1_UPPER = MDW0_UPPER + MASTER1_DATA_WIDTH;
  localparam [12:0] MDW2_UPPER = MDW1_UPPER + MASTER2_DATA_WIDTH;
  localparam [12:0] MDW3_UPPER = MDW2_UPPER + MASTER3_DATA_WIDTH;
  localparam [12:0] MDW4_UPPER = MDW3_UPPER + MASTER4_DATA_WIDTH;  
  localparam [12:0] MDW5_UPPER = MDW4_UPPER + MASTER5_DATA_WIDTH;
  localparam [12:0] MDW6_UPPER = MDW5_UPPER + MASTER6_DATA_WIDTH;
  localparam [12:0] MDW7_UPPER = MDW6_UPPER + MASTER7_DATA_WIDTH;

  localparam integer SLAVE_DATA_WIDTH_PORT = ( SLAVE31_DATA_WIDTH + SLAVE30_DATA_WIDTH + SLAVE29_DATA_WIDTH + SLAVE28_DATA_WIDTH + SLAVE27_DATA_WIDTH +
                                               SLAVE26_DATA_WIDTH + SLAVE25_DATA_WIDTH + SLAVE24_DATA_WIDTH + SLAVE23_DATA_WIDTH + SLAVE22_DATA_WIDTH +
                                               SLAVE21_DATA_WIDTH + SLAVE20_DATA_WIDTH + SLAVE19_DATA_WIDTH + SLAVE18_DATA_WIDTH + SLAVE17_DATA_WIDTH +
                                               SLAVE16_DATA_WIDTH + SLAVE15_DATA_WIDTH + SLAVE14_DATA_WIDTH + SLAVE13_DATA_WIDTH + SLAVE12_DATA_WIDTH +
                                               SLAVE11_DATA_WIDTH + SLAVE10_DATA_WIDTH + SLAVE9_DATA_WIDTH + SLAVE8_DATA_WIDTH +
                                               SLAVE7_DATA_WIDTH + SLAVE6_DATA_WIDTH + SLAVE5_DATA_WIDTH + SLAVE4_DATA_WIDTH +
                                               SLAVE3_DATA_WIDTH + SLAVE2_DATA_WIDTH + SLAVE1_DATA_WIDTH + SLAVE0_DATA_WIDTH);
  
  localparam [12:0] SDW0_UPPER = SLAVE0_DATA_WIDTH;
  localparam [12:0] SDW1_UPPER = SDW0_UPPER + SLAVE1_DATA_WIDTH;
  localparam [12:0] SDW2_UPPER = SDW1_UPPER + SLAVE2_DATA_WIDTH;
  localparam [12:0] SDW3_UPPER = SDW2_UPPER + SLAVE3_DATA_WIDTH;
  localparam [12:0] SDW4_UPPER = SDW3_UPPER + SLAVE4_DATA_WIDTH;
  localparam [12:0] SDW5_UPPER = SDW4_UPPER + SLAVE5_DATA_WIDTH;
  localparam [12:0] SDW6_UPPER = SDW5_UPPER + SLAVE6_DATA_WIDTH;
  localparam [12:0] SDW7_UPPER = SDW6_UPPER + SLAVE7_DATA_WIDTH;

  localparam [12:0] SDW8_UPPER  = SDW7_UPPER  + SLAVE8_DATA_WIDTH;
  localparam [12:0] SDW9_UPPER  = SDW8_UPPER  + SLAVE9_DATA_WIDTH;
  localparam [12:0] SDW10_UPPER = SDW9_UPPER  + SLAVE10_DATA_WIDTH;
  localparam [12:0] SDW11_UPPER = SDW10_UPPER + SLAVE11_DATA_WIDTH;
  localparam [12:0] SDW12_UPPER = SDW11_UPPER + SLAVE12_DATA_WIDTH;
  localparam [12:0] SDW13_UPPER = SDW12_UPPER + SLAVE13_DATA_WIDTH;
  localparam [12:0] SDW14_UPPER = SDW13_UPPER + SLAVE14_DATA_WIDTH;
  localparam [12:0] SDW15_UPPER = SDW14_UPPER + SLAVE15_DATA_WIDTH;
  localparam [12:0] SDW16_UPPER = SDW15_UPPER + SLAVE16_DATA_WIDTH;
  localparam [12:0] SDW17_UPPER = SDW16_UPPER + SLAVE17_DATA_WIDTH;
  localparam [12:0] SDW18_UPPER = SDW17_UPPER + SLAVE18_DATA_WIDTH;
  localparam [12:0] SDW19_UPPER = SDW18_UPPER + SLAVE19_DATA_WIDTH;
  localparam [12:0] SDW20_UPPER = SDW19_UPPER + SLAVE20_DATA_WIDTH;
  localparam [12:0] SDW21_UPPER = SDW20_UPPER + SLAVE21_DATA_WIDTH;
  localparam [12:0] SDW22_UPPER = SDW21_UPPER + SLAVE22_DATA_WIDTH;
  localparam [12:0] SDW23_UPPER = SDW22_UPPER + SLAVE23_DATA_WIDTH;
  localparam [12:0] SDW24_UPPER = SDW23_UPPER + SLAVE24_DATA_WIDTH;
  localparam [12:0] SDW25_UPPER = SDW24_UPPER + SLAVE25_DATA_WIDTH;
  localparam [12:0] SDW26_UPPER = SDW25_UPPER + SLAVE26_DATA_WIDTH;
  localparam [12:0] SDW27_UPPER = SDW26_UPPER + SLAVE27_DATA_WIDTH;
  localparam [12:0] SDW28_UPPER = SDW27_UPPER + SLAVE28_DATA_WIDTH;
  localparam [12:0] SDW29_UPPER = SDW28_UPPER + SLAVE29_DATA_WIDTH;
  localparam [12:0] SDW30_UPPER = SDW29_UPPER + SLAVE30_DATA_WIDTH;
  localparam [12:0] SDW31_UPPER = SDW30_UPPER + SLAVE31_DATA_WIDTH;

  localparam [13*NUM_MASTERS-1:0] MDW_UPPER_VEC = { MDW7_UPPER, MDW6_UPPER, MDW5_UPPER, MDW4_UPPER, MDW3_UPPER, MDW2_UPPER, MDW1_UPPER, MDW0_UPPER };
  localparam [13*NUM_MASTERS-1:0] MDW_LOWER_VEC = { MDW6_UPPER, MDW5_UPPER, MDW4_UPPER, MDW3_UPPER, MDW2_UPPER, MDW1_UPPER, MDW0_UPPER, 13'h0 };
  
  localparam [13*NUM_SLAVES-1:0] SDW_UPPER_VEC = { SDW31_UPPER, SDW30_UPPER, SDW29_UPPER, SDW28_UPPER, 
                                          SDW27_UPPER, SDW26_UPPER, SDW25_UPPER, SDW24_UPPER, 
                                          SDW23_UPPER, SDW22_UPPER, SDW21_UPPER, SDW20_UPPER,
                                          SDW19_UPPER, SDW18_UPPER, SDW17_UPPER, SDW16_UPPER, 
                                          SDW15_UPPER, SDW14_UPPER, SDW13_UPPER, SDW12_UPPER, 
                                          SDW11_UPPER, SDW10_UPPER, SDW9_UPPER, SDW8_UPPER, 
                                          SDW7_UPPER, SDW6_UPPER, SDW5_UPPER, SDW4_UPPER, 
                                          SDW3_UPPER, SDW2_UPPER, SDW1_UPPER, SDW0_UPPER  };
                                          
  localparam [13*NUM_SLAVES-1:0] SDW_LOWER_VEC = { SDW30_UPPER, SDW29_UPPER, SDW28_UPPER, SDW27_UPPER, 
                                          SDW26_UPPER, SDW25_UPPER, SDW24_UPPER, SDW23_UPPER, 
                                          SDW22_UPPER, SDW21_UPPER, SDW20_UPPER, SDW19_UPPER, 
                                          SDW18_UPPER, SDW17_UPPER, SDW16_UPPER, SDW15_UPPER, 
                                          SDW14_UPPER, SDW13_UPPER, SDW12_UPPER, SDW11_UPPER, 
                                          SDW10_UPPER, SDW9_UPPER, SDW8_UPPER, SDW7_UPPER, 
                                          SDW6_UPPER, SDW5_UPPER, SDW4_UPPER,SDW3_UPPER, 
                                          SDW2_UPPER, SDW1_UPPER, SDW0_UPPER, 13'h0 };
  
  localparam integer MASTER_STRB_WIDTH_PORT = ( MASTER0_DATA_WIDTH/8 + MASTER1_DATA_WIDTH/8 + MASTER2_DATA_WIDTH/8 + MASTER3_DATA_WIDTH/8 + MASTER4_DATA_WIDTH/8 + MASTER5_DATA_WIDTH/8 + MASTER6_DATA_WIDTH/8 + MASTER7_DATA_WIDTH/8);
  
  localparam integer SLAVE_STRB_WIDTH_PORT = ( SLAVE31_DATA_WIDTH/8 + SLAVE30_DATA_WIDTH/8 + SLAVE29_DATA_WIDTH/8 + SLAVE28_DATA_WIDTH/8 + 
                                               SLAVE27_DATA_WIDTH/8 + SLAVE26_DATA_WIDTH/8 + SLAVE25_DATA_WIDTH/8 + SLAVE24_DATA_WIDTH/8 + 
                                               SLAVE23_DATA_WIDTH/8 + SLAVE22_DATA_WIDTH/8 + SLAVE21_DATA_WIDTH/8 + SLAVE20_DATA_WIDTH/8 + 
                                               SLAVE19_DATA_WIDTH/8 + SLAVE18_DATA_WIDTH/8 + SLAVE17_DATA_WIDTH/8 + SLAVE16_DATA_WIDTH/8 + 
                                               SLAVE15_DATA_WIDTH/8 + SLAVE14_DATA_WIDTH/8 + SLAVE13_DATA_WIDTH/8 + SLAVE12_DATA_WIDTH/8 + 
                                               SLAVE11_DATA_WIDTH/8 + SLAVE10_DATA_WIDTH/8 + SLAVE9_DATA_WIDTH/8 + SLAVE8_DATA_WIDTH/8 + 
                                               SLAVE7_DATA_WIDTH/8 + SLAVE6_DATA_WIDTH/8 + SLAVE5_DATA_WIDTH/8 + SLAVE4_DATA_WIDTH/8 + 
                                               SLAVE3_DATA_WIDTH/8 + SLAVE2_DATA_WIDTH/8 + SLAVE1_DATA_WIDTH/8 + SLAVE0_DATA_WIDTH/8 );

  localparam [NUM_SLAVES-1:0]   MASTER0_WRITE_CONNECTIVITY   = { MASTER0_WRITE_SLAVE31, MASTER0_WRITE_SLAVE30, MASTER0_WRITE_SLAVE29, MASTER0_WRITE_SLAVE28, MASTER0_WRITE_SLAVE27, MASTER0_WRITE_SLAVE26, MASTER0_WRITE_SLAVE25, MASTER0_WRITE_SLAVE24, 
                                                                 MASTER0_WRITE_SLAVE23, MASTER0_WRITE_SLAVE22, MASTER0_WRITE_SLAVE21, MASTER0_WRITE_SLAVE20, MASTER0_WRITE_SLAVE19, MASTER0_WRITE_SLAVE18, MASTER0_WRITE_SLAVE17, MASTER0_WRITE_SLAVE16, 
                                                                 MASTER0_WRITE_SLAVE15, MASTER0_WRITE_SLAVE14, MASTER0_WRITE_SLAVE13, MASTER0_WRITE_SLAVE12, MASTER0_WRITE_SLAVE11, MASTER0_WRITE_SLAVE10, MASTER0_WRITE_SLAVE9,  MASTER0_WRITE_SLAVE8,  
                                                                 MASTER0_WRITE_SLAVE7,  MASTER0_WRITE_SLAVE6,  MASTER0_WRITE_SLAVE5,  MASTER0_WRITE_SLAVE4,  MASTER0_WRITE_SLAVE3,  MASTER0_WRITE_SLAVE2,  MASTER0_WRITE_SLAVE1,  MASTER0_WRITE_SLAVE0 } ;

  localparam [NUM_SLAVES-1:0]   MASTER1_WRITE_CONNECTIVITY   = { MASTER1_WRITE_SLAVE31, MASTER1_WRITE_SLAVE30, MASTER1_WRITE_SLAVE29, MASTER1_WRITE_SLAVE28, MASTER1_WRITE_SLAVE27, MASTER1_WRITE_SLAVE26, MASTER1_WRITE_SLAVE25, MASTER1_WRITE_SLAVE24, 
                                                                 MASTER1_WRITE_SLAVE23, MASTER1_WRITE_SLAVE22, MASTER1_WRITE_SLAVE21, MASTER1_WRITE_SLAVE20, MASTER1_WRITE_SLAVE19, MASTER1_WRITE_SLAVE18, MASTER1_WRITE_SLAVE17, MASTER1_WRITE_SLAVE16, 
                                                                 MASTER1_WRITE_SLAVE15, MASTER1_WRITE_SLAVE14, MASTER1_WRITE_SLAVE13, MASTER1_WRITE_SLAVE12, MASTER1_WRITE_SLAVE11, MASTER1_WRITE_SLAVE10, MASTER1_WRITE_SLAVE9,  MASTER1_WRITE_SLAVE8,  
                                                                 MASTER1_WRITE_SLAVE7,  MASTER1_WRITE_SLAVE6,  MASTER1_WRITE_SLAVE5,  MASTER1_WRITE_SLAVE4,  MASTER1_WRITE_SLAVE3,  MASTER1_WRITE_SLAVE2,  MASTER1_WRITE_SLAVE1,  MASTER1_WRITE_SLAVE0 };
  
  localparam [NUM_SLAVES-1:0]   MASTER2_WRITE_CONNECTIVITY   = { MASTER2_WRITE_SLAVE31, MASTER2_WRITE_SLAVE30, MASTER2_WRITE_SLAVE29, MASTER2_WRITE_SLAVE28, MASTER2_WRITE_SLAVE27, MASTER2_WRITE_SLAVE26, MASTER2_WRITE_SLAVE25, MASTER2_WRITE_SLAVE24, 
                                                                 MASTER2_WRITE_SLAVE23, MASTER2_WRITE_SLAVE22, MASTER2_WRITE_SLAVE21, MASTER2_WRITE_SLAVE20, MASTER2_WRITE_SLAVE19, MASTER2_WRITE_SLAVE18, MASTER2_WRITE_SLAVE17, MASTER2_WRITE_SLAVE16, 
                                                                 MASTER2_WRITE_SLAVE15, MASTER2_WRITE_SLAVE14, MASTER2_WRITE_SLAVE13, MASTER2_WRITE_SLAVE12, MASTER2_WRITE_SLAVE11, MASTER2_WRITE_SLAVE10, MASTER2_WRITE_SLAVE9,  MASTER2_WRITE_SLAVE8,  
                                                                 MASTER2_WRITE_SLAVE7,  MASTER2_WRITE_SLAVE6,  MASTER2_WRITE_SLAVE5,  MASTER2_WRITE_SLAVE4,  MASTER2_WRITE_SLAVE3,  MASTER2_WRITE_SLAVE2,  MASTER2_WRITE_SLAVE1,  MASTER2_WRITE_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER3_WRITE_CONNECTIVITY   = { MASTER3_WRITE_SLAVE31, MASTER3_WRITE_SLAVE30, MASTER3_WRITE_SLAVE29, MASTER3_WRITE_SLAVE28, MASTER3_WRITE_SLAVE27, MASTER3_WRITE_SLAVE26, MASTER3_WRITE_SLAVE25, MASTER3_WRITE_SLAVE24, 
                                                                 MASTER3_WRITE_SLAVE23, MASTER3_WRITE_SLAVE22, MASTER3_WRITE_SLAVE21, MASTER3_WRITE_SLAVE20, MASTER3_WRITE_SLAVE19, MASTER3_WRITE_SLAVE18, MASTER3_WRITE_SLAVE17, MASTER3_WRITE_SLAVE16, 
                                                                 MASTER3_WRITE_SLAVE15, MASTER3_WRITE_SLAVE14, MASTER3_WRITE_SLAVE13, MASTER3_WRITE_SLAVE12, MASTER3_WRITE_SLAVE11, MASTER3_WRITE_SLAVE10, MASTER3_WRITE_SLAVE9,  MASTER3_WRITE_SLAVE8,  
                                                                 MASTER3_WRITE_SLAVE7,  MASTER3_WRITE_SLAVE6,  MASTER3_WRITE_SLAVE5,  MASTER3_WRITE_SLAVE4,  MASTER3_WRITE_SLAVE3,  MASTER3_WRITE_SLAVE2,  MASTER3_WRITE_SLAVE1,  MASTER3_WRITE_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER4_WRITE_CONNECTIVITY   = { MASTER4_WRITE_SLAVE31, MASTER4_WRITE_SLAVE30, MASTER4_WRITE_SLAVE29, MASTER4_WRITE_SLAVE28, MASTER4_WRITE_SLAVE27, MASTER4_WRITE_SLAVE26, MASTER4_WRITE_SLAVE25, MASTER4_WRITE_SLAVE24, 
                                                                 MASTER4_WRITE_SLAVE23, MASTER4_WRITE_SLAVE22, MASTER4_WRITE_SLAVE21, MASTER4_WRITE_SLAVE20, MASTER4_WRITE_SLAVE19, MASTER4_WRITE_SLAVE18, MASTER4_WRITE_SLAVE17, MASTER4_WRITE_SLAVE16, 
                                                                 MASTER4_WRITE_SLAVE15, MASTER4_WRITE_SLAVE14, MASTER4_WRITE_SLAVE13, MASTER4_WRITE_SLAVE12, MASTER4_WRITE_SLAVE11, MASTER4_WRITE_SLAVE10, MASTER4_WRITE_SLAVE9,  MASTER4_WRITE_SLAVE8,  
                                                                 MASTER4_WRITE_SLAVE7,  MASTER4_WRITE_SLAVE6,  MASTER4_WRITE_SLAVE5,  MASTER4_WRITE_SLAVE4,  MASTER4_WRITE_SLAVE3,  MASTER4_WRITE_SLAVE2,  MASTER4_WRITE_SLAVE1,  MASTER4_WRITE_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER5_WRITE_CONNECTIVITY   = { MASTER5_WRITE_SLAVE31, MASTER5_WRITE_SLAVE30, MASTER5_WRITE_SLAVE29, MASTER5_WRITE_SLAVE28, MASTER5_WRITE_SLAVE27, MASTER5_WRITE_SLAVE26, MASTER5_WRITE_SLAVE25, MASTER5_WRITE_SLAVE24, 
                                                                 MASTER5_WRITE_SLAVE23, MASTER5_WRITE_SLAVE22, MASTER5_WRITE_SLAVE21, MASTER5_WRITE_SLAVE20, MASTER5_WRITE_SLAVE19, MASTER5_WRITE_SLAVE18, MASTER5_WRITE_SLAVE17, MASTER5_WRITE_SLAVE16, 
                                                                 MASTER5_WRITE_SLAVE15, MASTER5_WRITE_SLAVE14, MASTER5_WRITE_SLAVE13, MASTER5_WRITE_SLAVE12, MASTER5_WRITE_SLAVE11, MASTER5_WRITE_SLAVE10, MASTER5_WRITE_SLAVE9,  MASTER5_WRITE_SLAVE8,  
                                                                 MASTER5_WRITE_SLAVE7,  MASTER5_WRITE_SLAVE6,  MASTER5_WRITE_SLAVE5,  MASTER5_WRITE_SLAVE4,  MASTER5_WRITE_SLAVE3,  MASTER5_WRITE_SLAVE2,  MASTER5_WRITE_SLAVE1,  MASTER5_WRITE_SLAVE0 };
                            
  localparam [NUM_SLAVES-1:0]   MASTER6_WRITE_CONNECTIVITY   = { MASTER6_WRITE_SLAVE31, MASTER6_WRITE_SLAVE30, MASTER6_WRITE_SLAVE29, MASTER6_WRITE_SLAVE28, MASTER6_WRITE_SLAVE27, MASTER6_WRITE_SLAVE26, MASTER6_WRITE_SLAVE25, MASTER6_WRITE_SLAVE24, 
                                                                 MASTER6_WRITE_SLAVE23, MASTER6_WRITE_SLAVE22, MASTER6_WRITE_SLAVE21, MASTER6_WRITE_SLAVE20, MASTER6_WRITE_SLAVE19, MASTER6_WRITE_SLAVE18, MASTER6_WRITE_SLAVE17, MASTER6_WRITE_SLAVE16, 
                                                                 MASTER6_WRITE_SLAVE15, MASTER6_WRITE_SLAVE14, MASTER6_WRITE_SLAVE13, MASTER6_WRITE_SLAVE12, MASTER6_WRITE_SLAVE11, MASTER6_WRITE_SLAVE10, MASTER6_WRITE_SLAVE9,  MASTER6_WRITE_SLAVE8,  
                                                                 MASTER6_WRITE_SLAVE7,  MASTER6_WRITE_SLAVE6,  MASTER6_WRITE_SLAVE5,  MASTER6_WRITE_SLAVE4,  MASTER6_WRITE_SLAVE3,  MASTER6_WRITE_SLAVE2,  MASTER6_WRITE_SLAVE1,  MASTER6_WRITE_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER7_WRITE_CONNECTIVITY   = { MASTER7_WRITE_SLAVE31, MASTER7_WRITE_SLAVE30, MASTER7_WRITE_SLAVE29, MASTER7_WRITE_SLAVE28, MASTER7_WRITE_SLAVE27, MASTER7_WRITE_SLAVE26, MASTER7_WRITE_SLAVE25, MASTER7_WRITE_SLAVE24, 
                                                                 MASTER7_WRITE_SLAVE23, MASTER7_WRITE_SLAVE22, MASTER7_WRITE_SLAVE21, MASTER7_WRITE_SLAVE20, MASTER7_WRITE_SLAVE19, MASTER7_WRITE_SLAVE18, MASTER7_WRITE_SLAVE17, MASTER7_WRITE_SLAVE16, 
                                                                 MASTER7_WRITE_SLAVE15, MASTER7_WRITE_SLAVE14, MASTER7_WRITE_SLAVE13, MASTER7_WRITE_SLAVE12, MASTER7_WRITE_SLAVE11, MASTER7_WRITE_SLAVE10, MASTER7_WRITE_SLAVE9,  MASTER7_WRITE_SLAVE8,  
                                                                 MASTER7_WRITE_SLAVE7,  MASTER7_WRITE_SLAVE6,  MASTER7_WRITE_SLAVE5,  MASTER7_WRITE_SLAVE4,  MASTER7_WRITE_SLAVE3,  MASTER7_WRITE_SLAVE2,  MASTER7_WRITE_SLAVE1,  MASTER7_WRITE_SLAVE0 };


  localparam [NUM_SLAVES-1:0]   MASTER0_READ_CONNECTIVITY   = { MASTER0_READ_SLAVE31, MASTER0_READ_SLAVE30, MASTER0_READ_SLAVE29, MASTER0_READ_SLAVE28, MASTER0_READ_SLAVE27, MASTER0_READ_SLAVE26, MASTER0_READ_SLAVE25, MASTER0_READ_SLAVE24, 
                                                                MASTER0_READ_SLAVE23, MASTER0_READ_SLAVE22, MASTER0_READ_SLAVE21, MASTER0_READ_SLAVE20, MASTER0_READ_SLAVE19, MASTER0_READ_SLAVE18, MASTER0_READ_SLAVE17, MASTER0_READ_SLAVE16, 
                                                                MASTER0_READ_SLAVE15, MASTER0_READ_SLAVE14, MASTER0_READ_SLAVE13, MASTER0_READ_SLAVE12, MASTER0_READ_SLAVE11, MASTER0_READ_SLAVE10, MASTER0_READ_SLAVE9,  MASTER0_READ_SLAVE8,  
                                                                MASTER0_READ_SLAVE7,  MASTER0_READ_SLAVE6,  MASTER0_READ_SLAVE5,  MASTER0_READ_SLAVE4,  MASTER0_READ_SLAVE3,  MASTER0_READ_SLAVE2,  MASTER0_READ_SLAVE1,  MASTER0_READ_SLAVE0 } ;

  localparam [NUM_SLAVES-1:0]   MASTER1_READ_CONNECTIVITY   = { MASTER1_READ_SLAVE31, MASTER1_READ_SLAVE30, MASTER1_READ_SLAVE29, MASTER1_READ_SLAVE28, MASTER1_READ_SLAVE27, MASTER1_READ_SLAVE26, MASTER1_READ_SLAVE25, MASTER1_READ_SLAVE24, 
                                                                MASTER1_READ_SLAVE23, MASTER1_READ_SLAVE22, MASTER1_READ_SLAVE21, MASTER1_READ_SLAVE20, MASTER1_READ_SLAVE19, MASTER1_READ_SLAVE18, MASTER1_READ_SLAVE17, MASTER1_READ_SLAVE16, 
                                                                MASTER1_READ_SLAVE15, MASTER1_READ_SLAVE14, MASTER1_READ_SLAVE13, MASTER1_READ_SLAVE12, MASTER1_READ_SLAVE11, MASTER1_READ_SLAVE10, MASTER1_READ_SLAVE9,  MASTER1_READ_SLAVE8,  
                                                                MASTER1_READ_SLAVE7,  MASTER1_READ_SLAVE6,  MASTER1_READ_SLAVE5,  MASTER1_READ_SLAVE4,  MASTER1_READ_SLAVE3,  MASTER1_READ_SLAVE2,  MASTER1_READ_SLAVE1,  MASTER1_READ_SLAVE0 };
  
  localparam [NUM_SLAVES-1:0]   MASTER2_READ_CONNECTIVITY   = { MASTER2_READ_SLAVE31, MASTER2_READ_SLAVE30, MASTER2_READ_SLAVE29, MASTER2_READ_SLAVE28, MASTER2_READ_SLAVE27, MASTER2_READ_SLAVE26, MASTER2_READ_SLAVE25, MASTER2_READ_SLAVE24, 
                                                                MASTER2_READ_SLAVE23, MASTER2_READ_SLAVE22, MASTER2_READ_SLAVE21, MASTER2_READ_SLAVE20, MASTER2_READ_SLAVE19, MASTER2_READ_SLAVE18, MASTER2_READ_SLAVE17, MASTER2_READ_SLAVE16, 
                                                                MASTER2_READ_SLAVE15, MASTER2_READ_SLAVE14, MASTER2_READ_SLAVE13, MASTER2_READ_SLAVE12, MASTER2_READ_SLAVE11, MASTER2_READ_SLAVE10, MASTER2_READ_SLAVE9,  MASTER2_READ_SLAVE8,  
                                                                MASTER2_READ_SLAVE7,  MASTER2_READ_SLAVE6,  MASTER2_READ_SLAVE5,  MASTER2_READ_SLAVE4,  MASTER2_READ_SLAVE3,  MASTER2_READ_SLAVE2,  MASTER2_READ_SLAVE1,  MASTER2_READ_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER3_READ_CONNECTIVITY   = { MASTER3_READ_SLAVE31, MASTER3_READ_SLAVE30, MASTER3_READ_SLAVE29, MASTER3_READ_SLAVE28, MASTER3_READ_SLAVE27, MASTER3_READ_SLAVE26, MASTER3_READ_SLAVE25, MASTER3_READ_SLAVE24, 
                                                                MASTER3_READ_SLAVE23, MASTER3_READ_SLAVE22, MASTER3_READ_SLAVE21, MASTER3_READ_SLAVE20, MASTER3_READ_SLAVE19, MASTER3_READ_SLAVE18, MASTER3_READ_SLAVE17, MASTER3_READ_SLAVE16, 
                                                                MASTER3_READ_SLAVE15, MASTER3_READ_SLAVE14, MASTER3_READ_SLAVE13, MASTER3_READ_SLAVE12, MASTER3_READ_SLAVE11, MASTER3_READ_SLAVE10, MASTER3_READ_SLAVE9,  MASTER3_READ_SLAVE8,  
                                                                MASTER3_READ_SLAVE7,  MASTER3_READ_SLAVE6,  MASTER3_READ_SLAVE5,  MASTER3_READ_SLAVE4,  MASTER3_READ_SLAVE3,  MASTER3_READ_SLAVE2,  MASTER3_READ_SLAVE1,  MASTER3_READ_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER4_READ_CONNECTIVITY   = { MASTER4_READ_SLAVE31, MASTER4_READ_SLAVE30, MASTER4_READ_SLAVE29, MASTER4_READ_SLAVE28, MASTER4_READ_SLAVE27, MASTER4_READ_SLAVE26, MASTER4_READ_SLAVE25, MASTER4_READ_SLAVE24, 
                                                                MASTER4_READ_SLAVE23, MASTER4_READ_SLAVE22, MASTER4_READ_SLAVE21, MASTER4_READ_SLAVE20, MASTER4_READ_SLAVE19, MASTER4_READ_SLAVE18, MASTER4_READ_SLAVE17, MASTER4_READ_SLAVE16, 
                                                                MASTER4_READ_SLAVE15, MASTER4_READ_SLAVE14, MASTER4_READ_SLAVE13, MASTER4_READ_SLAVE12, MASTER4_READ_SLAVE11, MASTER4_READ_SLAVE10, MASTER4_READ_SLAVE9,  MASTER4_READ_SLAVE8,  
                                                                MASTER4_READ_SLAVE7,  MASTER4_READ_SLAVE6,  MASTER4_READ_SLAVE5,  MASTER4_READ_SLAVE4,  MASTER4_READ_SLAVE3,  MASTER4_READ_SLAVE2,  MASTER4_READ_SLAVE1,  MASTER4_READ_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER5_READ_CONNECTIVITY   = { MASTER5_READ_SLAVE31, MASTER5_READ_SLAVE30, MASTER5_READ_SLAVE29, MASTER5_READ_SLAVE28, MASTER5_READ_SLAVE27, MASTER5_READ_SLAVE26, MASTER5_READ_SLAVE25, MASTER5_READ_SLAVE24, 
                                                                MASTER5_READ_SLAVE23, MASTER5_READ_SLAVE22, MASTER5_READ_SLAVE21, MASTER5_READ_SLAVE20, MASTER5_READ_SLAVE19, MASTER5_READ_SLAVE18, MASTER5_READ_SLAVE17, MASTER5_READ_SLAVE16, 
                                                                MASTER5_READ_SLAVE15, MASTER5_READ_SLAVE14, MASTER5_READ_SLAVE13, MASTER5_READ_SLAVE12, MASTER5_READ_SLAVE11, MASTER5_READ_SLAVE10, MASTER5_READ_SLAVE9,  MASTER5_READ_SLAVE8,  
                                                                MASTER5_READ_SLAVE7,  MASTER5_READ_SLAVE6,  MASTER5_READ_SLAVE5,  MASTER5_READ_SLAVE4,  MASTER5_READ_SLAVE3,  MASTER5_READ_SLAVE2,  MASTER5_READ_SLAVE1,  MASTER5_READ_SLAVE0 };
                            
  localparam [NUM_SLAVES-1:0]   MASTER6_READ_CONNECTIVITY   = { MASTER6_READ_SLAVE31, MASTER6_READ_SLAVE30, MASTER6_READ_SLAVE29, MASTER6_READ_SLAVE28, MASTER6_READ_SLAVE27, MASTER6_READ_SLAVE26, MASTER6_READ_SLAVE25, MASTER6_READ_SLAVE24, 
                                                                MASTER6_READ_SLAVE23, MASTER6_READ_SLAVE22, MASTER6_READ_SLAVE21, MASTER6_READ_SLAVE20, MASTER6_READ_SLAVE19, MASTER6_READ_SLAVE18, MASTER6_READ_SLAVE17, MASTER6_READ_SLAVE16, 
                                                                MASTER6_READ_SLAVE15, MASTER6_READ_SLAVE14, MASTER6_READ_SLAVE13, MASTER6_READ_SLAVE12, MASTER6_READ_SLAVE11, MASTER6_READ_SLAVE10, MASTER6_READ_SLAVE9,  MASTER6_READ_SLAVE8,  
                                                                MASTER6_READ_SLAVE7,  MASTER6_READ_SLAVE6,  MASTER6_READ_SLAVE5,  MASTER6_READ_SLAVE4,  MASTER6_READ_SLAVE3,  MASTER6_READ_SLAVE2,  MASTER6_READ_SLAVE1,  MASTER6_READ_SLAVE0 };

  localparam [NUM_SLAVES-1:0]   MASTER7_READ_CONNECTIVITY   = { MASTER7_READ_SLAVE31, MASTER7_READ_SLAVE30, MASTER7_READ_SLAVE29, MASTER7_READ_SLAVE28, MASTER7_READ_SLAVE27, MASTER7_READ_SLAVE26, MASTER7_READ_SLAVE25, MASTER7_READ_SLAVE24, 
                                                                MASTER7_READ_SLAVE23, MASTER7_READ_SLAVE22, MASTER7_READ_SLAVE21, MASTER7_READ_SLAVE20, MASTER7_READ_SLAVE19, MASTER7_READ_SLAVE18, MASTER7_READ_SLAVE17, MASTER7_READ_SLAVE16, 
                                                                MASTER7_READ_SLAVE15, MASTER7_READ_SLAVE14, MASTER7_READ_SLAVE13, MASTER7_READ_SLAVE12, MASTER7_READ_SLAVE11, MASTER7_READ_SLAVE10, MASTER7_READ_SLAVE9,  MASTER7_READ_SLAVE8,  
                                                                MASTER7_READ_SLAVE7,  MASTER7_READ_SLAVE6,  MASTER7_READ_SLAVE5,  MASTER7_READ_SLAVE4,  MASTER7_READ_SLAVE3,  MASTER7_READ_SLAVE2,  MASTER7_READ_SLAVE1,  MASTER7_READ_SLAVE0 };
                            
  
  localparam [NUM_MASTERS*NUM_SLAVES-1:0] MASTER_WRITE_CONNECTIVITY = {  MASTER7_WRITE_CONNECTIVITY, MASTER6_WRITE_CONNECTIVITY, MASTER5_WRITE_CONNECTIVITY, MASTER4_WRITE_CONNECTIVITY, 
                                  MASTER3_WRITE_CONNECTIVITY, MASTER2_WRITE_CONNECTIVITY, MASTER1_WRITE_CONNECTIVITY, MASTER0_WRITE_CONNECTIVITY };  // bit per port indicating if a master can write to a slave port

  localparam [NUM_MASTERS*NUM_SLAVES-1:0] MASTER_READ_CONNECTIVITY  = {  MASTER7_READ_CONNECTIVITY, MASTER6_READ_CONNECTIVITY, MASTER5_READ_CONNECTIVITY, MASTER4_READ_CONNECTIVITY, 
                                  MASTER3_READ_CONNECTIVITY, MASTER2_READ_CONNECTIVITY, MASTER1_READ_CONNECTIVITY, MASTER0_READ_CONNECTIVITY };  // bit per port indicating if a master can write to a slave port

  localparam [NUM_MASTERS*8-1:0] MASTER_DEF_BURST_LEN = {    MASTER7_DEF_BURST_LEN,
                                      MASTER6_DEF_BURST_LEN,
                                      MASTER5_DEF_BURST_LEN,
                                      MASTER4_DEF_BURST_LEN,
                                      MASTER3_DEF_BURST_LEN,
                                      MASTER2_DEF_BURST_LEN,
                                      MASTER1_DEF_BURST_LEN,
                                      MASTER0_DEF_BURST_LEN
                                    };


  localparam [NUM_SLAVES*14-1:0] SLAVE_DWC_DATA_FIFO_DEPTH = {  SLAVE31_DWC_DATA_FIFO_DEPTH, SLAVE30_DWC_DATA_FIFO_DEPTH, SLAVE29_DWC_DATA_FIFO_DEPTH, SLAVE28_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE27_DWC_DATA_FIFO_DEPTH, SLAVE26_DWC_DATA_FIFO_DEPTH, SLAVE25_DWC_DATA_FIFO_DEPTH, SLAVE24_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE23_DWC_DATA_FIFO_DEPTH, SLAVE22_DWC_DATA_FIFO_DEPTH, SLAVE21_DWC_DATA_FIFO_DEPTH, SLAVE20_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE19_DWC_DATA_FIFO_DEPTH, SLAVE18_DWC_DATA_FIFO_DEPTH, SLAVE17_DWC_DATA_FIFO_DEPTH, SLAVE16_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE15_DWC_DATA_FIFO_DEPTH, SLAVE14_DWC_DATA_FIFO_DEPTH, SLAVE13_DWC_DATA_FIFO_DEPTH, SLAVE12_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE11_DWC_DATA_FIFO_DEPTH, SLAVE10_DWC_DATA_FIFO_DEPTH, SLAVE9_DWC_DATA_FIFO_DEPTH, SLAVE8_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE7_DWC_DATA_FIFO_DEPTH, SLAVE6_DWC_DATA_FIFO_DEPTH, SLAVE5_DWC_DATA_FIFO_DEPTH, SLAVE4_DWC_DATA_FIFO_DEPTH, 
                                                                SLAVE3_DWC_DATA_FIFO_DEPTH, SLAVE2_DWC_DATA_FIFO_DEPTH, SLAVE1_DWC_DATA_FIFO_DEPTH, SLAVE0_DWC_DATA_FIFO_DEPTH
                                                               };

  localparam [NUM_MASTERS*14-1:0] MASTER_DWC_DATA_FIFO_DEPTH = {  MASTER7_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER6_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER5_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER4_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER3_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER2_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER1_DWC_DATA_FIFO_DEPTH,
                                                                  MASTER0_DWC_DATA_FIFO_DEPTH
                                                                  };

  localparam [NUM_SLAVES-1:0] S_CDC = { SLAVE31_CLOCK_DOMAIN_CROSSING,SLAVE30_CLOCK_DOMAIN_CROSSING, SLAVE29_CLOCK_DOMAIN_CROSSING, SLAVE28_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE27_CLOCK_DOMAIN_CROSSING, SLAVE26_CLOCK_DOMAIN_CROSSING, SLAVE25_CLOCK_DOMAIN_CROSSING, SLAVE24_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE23_CLOCK_DOMAIN_CROSSING, SLAVE22_CLOCK_DOMAIN_CROSSING, SLAVE21_CLOCK_DOMAIN_CROSSING, SLAVE20_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE19_CLOCK_DOMAIN_CROSSING, SLAVE18_CLOCK_DOMAIN_CROSSING, SLAVE17_CLOCK_DOMAIN_CROSSING, SLAVE16_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE15_CLOCK_DOMAIN_CROSSING, SLAVE14_CLOCK_DOMAIN_CROSSING, SLAVE13_CLOCK_DOMAIN_CROSSING, SLAVE12_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE11_CLOCK_DOMAIN_CROSSING, SLAVE10_CLOCK_DOMAIN_CROSSING, SLAVE9_CLOCK_DOMAIN_CROSSING, SLAVE8_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE7_CLOCK_DOMAIN_CROSSING, SLAVE6_CLOCK_DOMAIN_CROSSING, SLAVE5_CLOCK_DOMAIN_CROSSING, SLAVE4_CLOCK_DOMAIN_CROSSING, 
                                        SLAVE3_CLOCK_DOMAIN_CROSSING, SLAVE2_CLOCK_DOMAIN_CROSSING, SLAVE1_CLOCK_DOMAIN_CROSSING, SLAVE0_CLOCK_DOMAIN_CROSSING 
                                      };

  localparam [NUM_MASTERS-1:0] M_CDC = {MASTER7_CLOCK_DOMAIN_CROSSING, MASTER6_CLOCK_DOMAIN_CROSSING, MASTER5_CLOCK_DOMAIN_CROSSING, MASTER4_CLOCK_DOMAIN_CROSSING, MASTER3_CLOCK_DOMAIN_CROSSING,  MASTER2_CLOCK_DOMAIN_CROSSING, MASTER1_CLOCK_DOMAIN_CROSSING, MASTER0_CLOCK_DOMAIN_CROSSING};


  //===================================================================================================================================

  //================================================= Global Signals  ==============================================//
  input  wire                                                        ACLK;
  input  wire                                                        ARESETN;      // active low reset synchronoise to RE AClk - asserted async.
   
  //================================================= Master Ports  ================================================//
  // AHB interface
  input wire  [31:0]  MASTER0_HADDR,     MASTER1_HADDR,     MASTER2_HADDR,     MASTER3_HADDR,     MASTER4_HADDR,     MASTER5_HADDR,     MASTER6_HADDR,     MASTER7_HADDR;
  input wire  [2:0]   MASTER0_HBURST,    MASTER1_HBURST,    MASTER2_HBURST,    MASTER3_HBURST,    MASTER4_HBURST,    MASTER5_HBURST,    MASTER6_HBURST,    MASTER7_HBURST;
  input wire          MASTER0_HMASTLOCK, MASTER1_HMASTLOCK, MASTER2_HMASTLOCK, MASTER3_HMASTLOCK, MASTER4_HMASTLOCK, MASTER5_HMASTLOCK, MASTER6_HMASTLOCK, MASTER7_HMASTLOCK;
  input wire  [6:0]   MASTER0_HPROT,     MASTER1_HPROT,     MASTER2_HPROT,     MASTER3_HPROT,     MASTER4_HPROT,     MASTER5_HPROT,     MASTER6_HPROT,     MASTER7_HPROT;
  input wire  [2:0]   MASTER0_HSIZE,     MASTER1_HSIZE,     MASTER2_HSIZE,     MASTER3_HSIZE,     MASTER4_HSIZE,     MASTER5_HSIZE,     MASTER6_HSIZE,     MASTER7_HSIZE;
  input wire          MASTER0_HNONSEC,   MASTER1_HNONSEC,   MASTER2_HNONSEC,   MASTER3_HNONSEC,   MASTER4_HNONSEC,   MASTER5_HNONSEC,   MASTER6_HNONSEC,   MASTER7_HNONSEC;
  input wire  [1:0]   MASTER0_HTRANS,    MASTER1_HTRANS,    MASTER2_HTRANS,    MASTER3_HTRANS,    MASTER4_HTRANS,    MASTER5_HTRANS,    MASTER6_HTRANS,    MASTER7_HTRANS;
  input wire          MASTER0_HWRITE,    MASTER1_HWRITE,    MASTER2_HWRITE,    MASTER3_HWRITE,    MASTER4_HWRITE,    MASTER5_HWRITE,    MASTER6_HWRITE,    MASTER7_HWRITE;
  output wire         MASTER0_HREADY,    MASTER1_HREADY,    MASTER2_HREADY,    MASTER3_HREADY,    MASTER4_HREADY,    MASTER5_HREADY,    MASTER6_HREADY,    MASTER7_HREADY;
  output wire         MASTER0_HRESP,     MASTER1_HRESP,     MASTER2_HRESP,     MASTER3_HRESP,     MASTER4_HRESP,     MASTER5_HRESP,     MASTER6_HRESP,     MASTER7_HRESP;
  // output wire         MASTER0_HEXOKAY,   MASTER1_HEXOKAY,   MASTER2_HEXOKAY,   MASTER3_HEXOKAY,   MASTER4_HEXOKAY,   MASTER5_HEXOKAY,   MASTER6_HEXOKAY,   MASTER7_HEXOKAY;
  input wire          MASTER0_HSEL,      MASTER1_HSEL,      MASTER2_HSEL,      MASTER3_HSEL,      MASTER4_HSEL,      MASTER5_HSEL,      MASTER6_HSEL,      MASTER7_HSEL;
  // input wire          MASTER0_HEXCL,     MASTER1_HEXCL,     MASTER2_HEXCL,     MASTER3_HEXCL,     MASTER4_HEXCL,     MASTER5_HEXCL,     MASTER6_HEXCL,     MASTER7_HEXCL;

  // AHB data ports
  input  wire [MASTER0_DATA_WIDTH-1:0]    MASTER0_HWDATA;  
  input  wire [MASTER1_DATA_WIDTH-1:0]    MASTER1_HWDATA;  
  input  wire [MASTER2_DATA_WIDTH-1:0]    MASTER2_HWDATA;  
  input  wire [MASTER3_DATA_WIDTH-1:0]    MASTER3_HWDATA;  
  input  wire [MASTER4_DATA_WIDTH-1:0]    MASTER4_HWDATA;  
  input  wire [MASTER5_DATA_WIDTH-1:0]    MASTER5_HWDATA;  
  input  wire [MASTER6_DATA_WIDTH-1:0]    MASTER6_HWDATA;  
  input  wire [MASTER7_DATA_WIDTH-1:0]    MASTER7_HWDATA;

  output  wire [MASTER0_DATA_WIDTH-1:0]    MASTER0_HRDATA;  
  output  wire [MASTER1_DATA_WIDTH-1:0]    MASTER1_HRDATA;  
  output  wire [MASTER2_DATA_WIDTH-1:0]    MASTER2_HRDATA;  
  output  wire [MASTER3_DATA_WIDTH-1:0]    MASTER3_HRDATA;  
  output  wire [MASTER4_DATA_WIDTH-1:0]    MASTER4_HRDATA;  
  output  wire [MASTER5_DATA_WIDTH-1:0]    MASTER5_HRDATA;  
  output  wire [MASTER6_DATA_WIDTH-1:0]    MASTER6_HRDATA;  
  output  wire [MASTER7_DATA_WIDTH-1:0]    MASTER7_HRDATA;


  // Master Write Address Ports                
  input  wire [ID_WIDTH-1:0]    MASTER0_AWID,     MASTER1_AWID,     MASTER2_AWID,     MASTER3_AWID,     MASTER4_AWID,     MASTER5_AWID,     MASTER6_AWID,     MASTER7_AWID;
  input  wire [ADDR_WIDTH-1:0]  MASTER0_AWADDR,   MASTER1_AWADDR,   MASTER2_AWADDR,   MASTER3_AWADDR,   MASTER4_AWADDR,   MASTER5_AWADDR,   MASTER6_AWADDR,   MASTER7_AWADDR;
  input  wire [7:0]             MASTER0_AWLEN,    MASTER1_AWLEN,    MASTER2_AWLEN,    MASTER3_AWLEN,    MASTER4_AWLEN,    MASTER5_AWLEN,    MASTER6_AWLEN,    MASTER7_AWLEN;
  input  wire [2:0]             MASTER0_AWSIZE,   MASTER1_AWSIZE,   MASTER2_AWSIZE,   MASTER3_AWSIZE,   MASTER4_AWSIZE,   MASTER5_AWSIZE,   MASTER6_AWSIZE,   MASTER7_AWSIZE;
  input  wire [1:0]             MASTER0_AWBURST,  MASTER1_AWBURST,  MASTER2_AWBURST,  MASTER3_AWBURST,  MASTER4_AWBURST,  MASTER5_AWBURST,  MASTER6_AWBURST,  MASTER7_AWBURST;
  input  wire [1:0]             MASTER0_AWLOCK,   MASTER1_AWLOCK,   MASTER2_AWLOCK,   MASTER3_AWLOCK,   MASTER4_AWLOCK,   MASTER5_AWLOCK,   MASTER6_AWLOCK,   MASTER7_AWLOCK;
  input  wire [3:0]             MASTER0_AWCACHE,  MASTER1_AWCACHE,  MASTER2_AWCACHE,  MASTER3_AWCACHE,  MASTER4_AWCACHE,  MASTER5_AWCACHE,  MASTER6_AWCACHE,  MASTER7_AWCACHE;
  input  wire [2:0]             MASTER0_AWPROT,   MASTER1_AWPROT,   MASTER2_AWPROT,   MASTER3_AWPROT,   MASTER4_AWPROT,   MASTER5_AWPROT,   MASTER6_AWPROT,   MASTER7_AWPROT;
  input  wire [3:0]             MASTER0_AWREGION, MASTER1_AWREGION, MASTER2_AWREGION, MASTER3_AWREGION, MASTER4_AWREGION, MASTER5_AWREGION, MASTER6_AWREGION, MASTER7_AWREGION;
  input  wire [3:0]             MASTER0_AWQOS,    MASTER1_AWQOS,    MASTER2_AWQOS,    MASTER3_AWQOS,    MASTER4_AWQOS,    MASTER5_AWQOS,    MASTER6_AWQOS,    MASTER7_AWQOS;
  input  wire [USER_WIDTH-1:0]  MASTER0_AWUSER,   MASTER1_AWUSER,   MASTER2_AWUSER,   MASTER3_AWUSER,   MASTER4_AWUSER,   MASTER5_AWUSER,   MASTER6_AWUSER,   MASTER7_AWUSER;
  input  wire                   MASTER0_AWVALID,  MASTER1_AWVALID,  MASTER2_AWVALID,  MASTER3_AWVALID,  MASTER4_AWVALID,  MASTER5_AWVALID,  MASTER6_AWVALID,  MASTER7_AWVALID;
  output wire                   MASTER0_AWREADY,  MASTER1_AWREADY,  MASTER2_AWREADY,  MASTER3_AWREADY,  MASTER4_AWREADY,  MASTER5_AWREADY,  MASTER6_AWREADY,  MASTER7_AWREADY;
  input wire                    M_CLK0,           M_CLK1,           M_CLK2,           M_CLK3,           M_CLK4,           M_CLK5,           M_CLK6,           M_CLK7;
  
  input wire                    S_CLK0,  S_CLK1,  S_CLK2,  S_CLK3,  S_CLK4,  S_CLK5,  S_CLK6,  S_CLK7, 
                                S_CLK8,  S_CLK9,  S_CLK10, S_CLK11, S_CLK12, S_CLK13, S_CLK14, S_CLK15, 
                                S_CLK16, S_CLK17, S_CLK18, S_CLK19, S_CLK20, S_CLK21, S_CLK22, S_CLK23, 
                                S_CLK24, S_CLK25, S_CLK26, S_CLK27, S_CLK28, S_CLK29, S_CLK30, S_CLK31;

  // Master Write Data Ports
  input  wire [MASTER0_DATA_WIDTH-1:0]    MASTER0_WDATA;  
  input  wire [MASTER1_DATA_WIDTH-1:0]    MASTER1_WDATA;  
  input  wire [MASTER2_DATA_WIDTH-1:0]    MASTER2_WDATA;  
  input  wire [MASTER3_DATA_WIDTH-1:0]    MASTER3_WDATA;  
  input  wire [MASTER4_DATA_WIDTH-1:0]    MASTER4_WDATA;  
  input  wire [MASTER5_DATA_WIDTH-1:0]    MASTER5_WDATA;  
  input  wire [MASTER6_DATA_WIDTH-1:0]    MASTER6_WDATA;  
  input  wire [MASTER7_DATA_WIDTH-1:0]    MASTER7_WDATA;
  input  wire [(MASTER0_DATA_WIDTH/8)-1:0]  MASTER0_WSTRB;  
  input  wire [(MASTER1_DATA_WIDTH/8)-1:0]  MASTER1_WSTRB;  
  input  wire [(MASTER2_DATA_WIDTH/8)-1:0]  MASTER2_WSTRB;  
  input  wire [(MASTER3_DATA_WIDTH/8)-1:0]  MASTER3_WSTRB;  
  input  wire [(MASTER4_DATA_WIDTH/8)-1:0]  MASTER4_WSTRB;  
  input  wire [(MASTER5_DATA_WIDTH/8)-1:0]  MASTER5_WSTRB;  
  input  wire [(MASTER6_DATA_WIDTH/8)-1:0]  MASTER6_WSTRB;  
  input  wire [(MASTER7_DATA_WIDTH/8)-1:0]  MASTER7_WSTRB;
  input  wire                    MASTER0_WLAST,   MASTER1_WLAST,  MASTER2_WLAST,  MASTER3_WLAST,  MASTER4_WLAST,  MASTER5_WLAST,  MASTER6_WLAST,  MASTER7_WLAST;
  input  wire [USER_WIDTH-1:0]   MASTER0_WUSER,   MASTER1_WUSER,  MASTER2_WUSER,  MASTER3_WUSER,  MASTER4_WUSER,  MASTER5_WUSER,  MASTER6_WUSER,  MASTER7_WUSER;
  input  wire                    MASTER0_WVALID,  MASTER1_WVALID, MASTER2_WVALID, MASTER3_WVALID, MASTER4_WVALID, MASTER5_WVALID, MASTER6_WVALID, MASTER7_WVALID;
  output wire                    MASTER0_WREADY,  MASTER1_WREADY, MASTER2_WREADY, MASTER3_WREADY, MASTER4_WREADY, MASTER5_WREADY, MASTER6_WREADY, MASTER7_WREADY;
                 
  // Master Write Response Ports                
  output wire [ID_WIDTH-1:0]     MASTER0_BID,    MASTER1_BID,    MASTER2_BID,    MASTER3_BID,    MASTER4_BID,    MASTER5_BID,    MASTER6_BID,    MASTER7_BID;
  output wire [1:0]              MASTER0_BRESP,  MASTER1_BRESP,  MASTER2_BRESP,  MASTER3_BRESP,  MASTER4_BRESP,  MASTER5_BRESP,  MASTER6_BRESP,  MASTER7_BRESP;
  output wire [USER_WIDTH-1:0]   MASTER0_BUSER,  MASTER1_BUSER,  MASTER2_BUSER,  MASTER3_BUSER,  MASTER4_BUSER,  MASTER5_BUSER,  MASTER6_BUSER,  MASTER7_BUSER;
  output wire                    MASTER0_BVALID, MASTER1_BVALID, MASTER2_BVALID, MASTER3_BVALID, MASTER4_BVALID, MASTER5_BVALID, MASTER6_BVALID, MASTER7_BVALID;
  input  wire                    MASTER0_BREADY, MASTER1_BREADY, MASTER2_BREADY, MASTER3_BREADY, MASTER4_BREADY, MASTER5_BREADY, MASTER6_BREADY, MASTER7_BREADY;
                
  // Master Read Address Ports                
  input  wire [ID_WIDTH-1:0]    MASTER0_ARID,     MASTER1_ARID,     MASTER2_ARID,     MASTER3_ARID,     MASTER4_ARID,     MASTER5_ARID,     MASTER6_ARID,     MASTER7_ARID;
  input  wire [ADDR_WIDTH-1:0]  MASTER0_ARADDR,   MASTER1_ARADDR,   MASTER2_ARADDR,   MASTER3_ARADDR,   MASTER4_ARADDR,   MASTER5_ARADDR,   MASTER6_ARADDR,   MASTER7_ARADDR;
  input  wire [7:0]             MASTER0_ARLEN,    MASTER1_ARLEN,    MASTER2_ARLEN,    MASTER3_ARLEN,    MASTER4_ARLEN,    MASTER5_ARLEN,    MASTER6_ARLEN,    MASTER7_ARLEN;
  input  wire [2:0]             MASTER0_ARSIZE,   MASTER1_ARSIZE,   MASTER2_ARSIZE,   MASTER3_ARSIZE,   MASTER4_ARSIZE,   MASTER5_ARSIZE,   MASTER6_ARSIZE,   MASTER7_ARSIZE;
  input  wire [1:0]             MASTER0_ARBURST,  MASTER1_ARBURST,  MASTER2_ARBURST,  MASTER3_ARBURST,  MASTER4_ARBURST,  MASTER5_ARBURST,  MASTER6_ARBURST,  MASTER7_ARBURST;
  input  wire [1:0]             MASTER0_ARLOCK,   MASTER1_ARLOCK,   MASTER2_ARLOCK,   MASTER3_ARLOCK,   MASTER4_ARLOCK,   MASTER5_ARLOCK,   MASTER6_ARLOCK,   MASTER7_ARLOCK;
  input  wire [3:0]             MASTER0_ARCACHE,  MASTER1_ARCACHE,  MASTER2_ARCACHE,  MASTER3_ARCACHE,  MASTER4_ARCACHE,  MASTER5_ARCACHE,  MASTER6_ARCACHE,  MASTER7_ARCACHE;
  input  wire [2:0]             MASTER0_ARPROT,   MASTER1_ARPROT,   MASTER2_ARPROT,   MASTER3_ARPROT,   MASTER4_ARPROT,   MASTER5_ARPROT,   MASTER6_ARPROT,   MASTER7_ARPROT;
  input  wire [3:0]             MASTER0_ARREGION, MASTER1_ARREGION, MASTER2_ARREGION, MASTER3_ARREGION, MASTER4_ARREGION, MASTER5_ARREGION, MASTER6_ARREGION, MASTER7_ARREGION;
  input  wire [3:0]             MASTER0_ARQOS,    MASTER1_ARQOS,    MASTER2_ARQOS,    MASTER3_ARQOS,    MASTER4_ARQOS,    MASTER5_ARQOS,    MASTER6_ARQOS,    MASTER7_ARQOS;
  input  wire [USER_WIDTH-1:0]  MASTER0_ARUSER,   MASTER1_ARUSER,   MASTER2_ARUSER,   MASTER3_ARUSER,   MASTER4_ARUSER,   MASTER5_ARUSER,   MASTER6_ARUSER,   MASTER7_ARUSER;
  input  wire                   MASTER0_ARVALID,  MASTER1_ARVALID,  MASTER2_ARVALID,  MASTER3_ARVALID,  MASTER4_ARVALID,  MASTER5_ARVALID,  MASTER6_ARVALID,  MASTER7_ARVALID;
  output wire                   MASTER0_ARREADY,  MASTER1_ARREADY,  MASTER2_ARREADY,  MASTER3_ARREADY,  MASTER4_ARREADY,  MASTER5_ARREADY,  MASTER6_ARREADY,  MASTER7_ARREADY;
                
  // Master Read Data Ports                
  output wire [ID_WIDTH-1:0]             MASTER0_RID,  MASTER1_RID,  MASTER2_RID,  MASTER3_RID,  MASTER4_RID,  MASTER5_RID,  MASTER6_RID,  MASTER7_RID;
  output wire [MASTER0_DATA_WIDTH-1:0]   MASTER0_RDATA;
  output wire [MASTER1_DATA_WIDTH-1:0]   MASTER1_RDATA;  
  output wire [MASTER2_DATA_WIDTH-1:0]   MASTER2_RDATA;  
  output wire [MASTER3_DATA_WIDTH-1:0]   MASTER3_RDATA;  
  output wire [MASTER4_DATA_WIDTH-1:0]   MASTER4_RDATA;  
  output wire [MASTER5_DATA_WIDTH-1:0]   MASTER5_RDATA;  
  output wire [MASTER6_DATA_WIDTH-1:0]   MASTER6_RDATA;  
  output wire [MASTER7_DATA_WIDTH-1:0]   MASTER7_RDATA;
  output wire [1:0]                      MASTER0_RRESP,  MASTER1_RRESP,  MASTER2_RRESP,  MASTER3_RRESP,  MASTER4_RRESP,  MASTER5_RRESP,  MASTER6_RRESP,  MASTER7_RRESP;
  output wire                            MASTER0_RLAST,  MASTER1_RLAST,  MASTER2_RLAST,  MASTER3_RLAST,  MASTER4_RLAST,  MASTER5_RLAST,  MASTER6_RLAST,  MASTER7_RLAST;
  output wire [USER_WIDTH-1:0]           MASTER0_RUSER,  MASTER1_RUSER,  MASTER2_RUSER,  MASTER3_RUSER,  MASTER4_RUSER,  MASTER5_RUSER,  MASTER6_RUSER,  MASTER7_RUSER;
  output wire                            MASTER0_RVALID, MASTER1_RVALID, MASTER2_RVALID, MASTER3_RVALID, MASTER4_RVALID, MASTER5_RVALID, MASTER6_RVALID, MASTER7_RVALID;
  input  wire                            MASTER0_RREADY, MASTER1_RREADY, MASTER2_RREADY, MASTER3_RREADY, MASTER4_RREADY, MASTER5_RREADY, MASTER6_RREADY, MASTER7_RREADY;
                   

  //================================================ Slave Ports  ======================================================================//
   
  // Slave Write Address Port - Slave ID is composed of Master Port ID concatenated with transaction ID
  output wire [(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]  SLAVE0_AWID,     SLAVE1_AWID,     SLAVE2_AWID,      SLAVE3_AWID,     SLAVE4_AWID,     SLAVE5_AWID,     SLAVE6_AWID,     SLAVE7_AWID,
                                                  SLAVE8_AWID,     SLAVE9_AWID,     SLAVE10_AWID,     SLAVE11_AWID,    SLAVE12_AWID,    SLAVE13_AWID,    SLAVE14_AWID,    SLAVE15_AWID,
                                                  SLAVE16_AWID,    SLAVE17_AWID,    SLAVE18_AWID,     SLAVE19_AWID,    SLAVE20_AWID,    SLAVE21_AWID,    SLAVE22_AWID,    SLAVE23_AWID,
                                                  SLAVE24_AWID,    SLAVE25_AWID,    SLAVE26_AWID,     SLAVE27_AWID,    SLAVE28_AWID,    SLAVE29_AWID,    SLAVE30_AWID,    SLAVE31_AWID;
                                                  
  output wire [ADDR_WIDTH-1:0]    SLAVE0_AWADDR,   SLAVE1_AWADDR,   SLAVE2_AWADDR,   SLAVE3_AWADDR,    SLAVE4_AWADDR,   SLAVE5_AWADDR,   SLAVE6_AWADDR,   SLAVE7_AWADDR,
                                  SLAVE8_AWADDR,   SLAVE9_AWADDR,   SLAVE10_AWADDR,  SLAVE11_AWADDR,   SLAVE12_AWADDR,  SLAVE13_AWADDR,  SLAVE14_AWADDR,  SLAVE15_AWADDR,
                                  SLAVE16_AWADDR,  SLAVE17_AWADDR,  SLAVE18_AWADDR,  SLAVE19_AWADDR,   SLAVE20_AWADDR,  SLAVE21_AWADDR,  SLAVE22_AWADDR,  SLAVE23_AWADDR,
                                  SLAVE24_AWADDR,  SLAVE25_AWADDR,  SLAVE26_AWADDR,  SLAVE27_AWADDR,   SLAVE28_AWADDR,  SLAVE29_AWADDR,  SLAVE30_AWADDR,  SLAVE31_AWADDR;
                                                  
  output wire [7:0]               SLAVE0_AWLEN,    SLAVE1_AWLEN,    SLAVE2_AWLEN,    SLAVE3_AWLEN,    SLAVE4_AWLEN,    SLAVE5_AWLEN,    SLAVE6_AWLEN,    SLAVE7_AWLEN,
                                  SLAVE8_AWLEN,    SLAVE9_AWLEN,    SLAVE10_AWLEN,   SLAVE11_AWLEN,   SLAVE12_AWLEN,   SLAVE13_AWLEN,   SLAVE14_AWLEN,   SLAVE15_AWLEN,
                                  SLAVE16_AWLEN,   SLAVE17_AWLEN,   SLAVE18_AWLEN,   SLAVE19_AWLEN,   SLAVE20_AWLEN,   SLAVE21_AWLEN,   SLAVE22_AWLEN,   SLAVE23_AWLEN,
                                  SLAVE24_AWLEN,   SLAVE25_AWLEN,   SLAVE26_AWLEN,   SLAVE27_AWLEN,   SLAVE28_AWLEN,   SLAVE29_AWLEN,   SLAVE30_AWLEN,   SLAVE31_AWLEN;
                                                  
  
  output wire [2:0]               SLAVE0_AWSIZE,   SLAVE1_AWSIZE,   SLAVE2_AWSIZE,   SLAVE3_AWSIZE,   SLAVE4_AWSIZE,   SLAVE5_AWSIZE,   SLAVE6_AWSIZE,   SLAVE7_AWSIZE,
                                  SLAVE8_AWSIZE,   SLAVE9_AWSIZE,   SLAVE10_AWSIZE,  SLAVE11_AWSIZE,  SLAVE12_AWSIZE,  SLAVE13_AWSIZE,  SLAVE14_AWSIZE,  SLAVE15_AWSIZE,
                                  SLAVE16_AWSIZE,  SLAVE17_AWSIZE,  SLAVE18_AWSIZE,  SLAVE19_AWSIZE,  SLAVE20_AWSIZE,  SLAVE21_AWSIZE,  SLAVE22_AWSIZE,  SLAVE23_AWSIZE,
                                  SLAVE24_AWSIZE,  SLAVE25_AWSIZE,  SLAVE26_AWSIZE,  SLAVE27_AWSIZE,  SLAVE28_AWSIZE,  SLAVE29_AWSIZE,  SLAVE30_AWSIZE,  SLAVE31_AWSIZE;


  output wire [1:0]               SLAVE0_AWBURST,  SLAVE1_AWBURST,  SLAVE2_AWBURST,   SLAVE3_AWBURST,  SLAVE4_AWBURST,  SLAVE5_AWBURST,  SLAVE6_AWBURST,   SLAVE7_AWBURST,
                                  SLAVE8_AWBURST,  SLAVE9_AWBURST,  SLAVE10_AWBURST,  SLAVE11_AWBURST, SLAVE12_AWBURST, SLAVE13_AWBURST, SLAVE14_AWBURST,  SLAVE15_AWBURST,
                                  SLAVE16_AWBURST, SLAVE17_AWBURST, SLAVE18_AWBURST,  SLAVE19_AWBURST, SLAVE20_AWBURST, SLAVE21_AWBURST, SLAVE22_AWBURST,  SLAVE23_AWBURST,
                                  SLAVE24_AWBURST, SLAVE25_AWBURST, SLAVE26_AWBURST,  SLAVE27_AWBURST, SLAVE28_AWBURST, SLAVE29_AWBURST, SLAVE30_AWBURST,  SLAVE31_AWBURST;

  
  output wire [1:0]               SLAVE0_AWLOCK,   SLAVE1_AWLOCK,   SLAVE2_AWLOCK,   SLAVE3_AWLOCK,   SLAVE4_AWLOCK,   SLAVE5_AWLOCK,   SLAVE6_AWLOCK,   SLAVE7_AWLOCK,
                                  SLAVE8_AWLOCK,   SLAVE9_AWLOCK,   SLAVE10_AWLOCK,  SLAVE11_AWLOCK,  SLAVE12_AWLOCK,  SLAVE13_AWLOCK,  SLAVE14_AWLOCK,  SLAVE15_AWLOCK,
                                  SLAVE16_AWLOCK,  SLAVE17_AWLOCK,  SLAVE18_AWLOCK,  SLAVE19_AWLOCK,  SLAVE20_AWLOCK,  SLAVE21_AWLOCK,  SLAVE22_AWLOCK,  SLAVE23_AWLOCK,
                                  SLAVE24_AWLOCK,  SLAVE25_AWLOCK,  SLAVE26_AWLOCK,  SLAVE27_AWLOCK,  SLAVE28_AWLOCK,  SLAVE29_AWLOCK,  SLAVE30_AWLOCK,  SLAVE31_AWLOCK;

  
  output wire [3:0]               SLAVE0_AWCACHE,   SLAVE1_AWCACHE,   SLAVE2_AWCACHE,   SLAVE3_AWCACHE,   SLAVE4_AWCACHE,   SLAVE5_AWCACHE,   SLAVE6_AWCACHE,   SLAVE7_AWCACHE,
                                  SLAVE8_AWCACHE,   SLAVE9_AWCACHE,   SLAVE10_AWCACHE,  SLAVE11_AWCACHE,  SLAVE12_AWCACHE,  SLAVE13_AWCACHE,  SLAVE14_AWCACHE,  SLAVE15_AWCACHE,
                                  SLAVE16_AWCACHE,  SLAVE17_AWCACHE,  SLAVE18_AWCACHE,  SLAVE19_AWCACHE,  SLAVE20_AWCACHE,  SLAVE21_AWCACHE,  SLAVE22_AWCACHE,  SLAVE23_AWCACHE,
                                  SLAVE24_AWCACHE,  SLAVE25_AWCACHE,  SLAVE26_AWCACHE,  SLAVE27_AWCACHE,  SLAVE28_AWCACHE,  SLAVE29_AWCACHE,  SLAVE30_AWCACHE,  SLAVE31_AWCACHE;

  output wire [2:0]               SLAVE0_AWPROT,   SLAVE1_AWPROT,   SLAVE2_AWPROT,   SLAVE3_AWPROT,   SLAVE4_AWPROT,   SLAVE5_AWPROT,   SLAVE6_AWPROT,   SLAVE7_AWPROT,
                                  SLAVE8_AWPROT,   SLAVE9_AWPROT,   SLAVE10_AWPROT,  SLAVE11_AWPROT,  SLAVE12_AWPROT,  SLAVE13_AWPROT,  SLAVE14_AWPROT,  SLAVE15_AWPROT,
                                  SLAVE16_AWPROT,  SLAVE17_AWPROT,  SLAVE18_AWPROT,  SLAVE19_AWPROT,  SLAVE20_AWPROT,  SLAVE21_AWPROT,  SLAVE22_AWPROT,  SLAVE23_AWPROT,
                                  SLAVE24_AWPROT,  SLAVE25_AWPROT,  SLAVE26_AWPROT,  SLAVE27_AWPROT,  SLAVE28_AWPROT,  SLAVE29_AWPROT,  SLAVE30_AWPROT,  SLAVE31_AWPROT;


  output wire [3:0]               SLAVE0_AWREGION,   SLAVE1_AWREGION,   SLAVE2_AWREGION,   SLAVE3_AWREGION,   SLAVE4_AWREGION,   SLAVE5_AWREGION,   SLAVE6_AWREGION,   SLAVE7_AWREGION,
                                  SLAVE8_AWREGION,   SLAVE9_AWREGION,   SLAVE10_AWREGION,  SLAVE11_AWREGION,  SLAVE12_AWREGION,  SLAVE13_AWREGION,  SLAVE14_AWREGION,  SLAVE15_AWREGION,
                                  SLAVE16_AWREGION,  SLAVE17_AWREGION,  SLAVE18_AWREGION,  SLAVE19_AWREGION,  SLAVE20_AWREGION,  SLAVE21_AWREGION,  SLAVE22_AWREGION,  SLAVE23_AWREGION,
                                  SLAVE24_AWREGION,  SLAVE25_AWREGION,  SLAVE26_AWREGION,  SLAVE27_AWREGION,  SLAVE28_AWREGION,  SLAVE29_AWREGION,  SLAVE30_AWREGION,  SLAVE31_AWREGION;

  output wire [3:0]               SLAVE0_AWQOS,   SLAVE1_AWQOS,  SLAVE2_AWQOS,   SLAVE3_AWQOS,  SLAVE4_AWQOS,   SLAVE5_AWQOS,   SLAVE6_AWQOS,   SLAVE7_AWQOS,
                                  SLAVE8_AWQOS,   SLAVE9_AWQOS,  SLAVE10_AWQOS,  SLAVE11_AWQOS, SLAVE12_AWQOS,  SLAVE13_AWQOS,  SLAVE14_AWQOS,  SLAVE15_AWQOS,
                                  SLAVE16_AWQOS,  SLAVE17_AWQOS, SLAVE18_AWQOS,  SLAVE19_AWQOS, SLAVE20_AWQOS,  SLAVE21_AWQOS,  SLAVE22_AWQOS,  SLAVE23_AWQOS,  
                                  SLAVE24_AWQOS,  SLAVE25_AWQOS, SLAVE26_AWQOS,  SLAVE27_AWQOS, SLAVE28_AWQOS,  SLAVE29_AWQOS,  SLAVE30_AWQOS,   SLAVE31_AWQOS;
                                  
                                  
  output wire [USER_WIDTH-1:0]    SLAVE0_AWUSER,   SLAVE1_AWUSER,   SLAVE2_AWUSER,   SLAVE3_AWUSER,   SLAVE4_AWUSER,   SLAVE5_AWUSER,   SLAVE6_AWUSER,   SLAVE7_AWUSER,
                                  SLAVE8_AWUSER,   SLAVE9_AWUSER,   SLAVE10_AWUSER,  SLAVE11_AWUSER,  SLAVE12_AWUSER,  SLAVE13_AWUSER,  SLAVE14_AWUSER,  SLAVE15_AWUSER,
                                  SLAVE16_AWUSER,  SLAVE17_AWUSER,  SLAVE18_AWUSER,  SLAVE19_AWUSER,  SLAVE20_AWUSER,  SLAVE21_AWUSER,  SLAVE22_AWUSER,  SLAVE23_AWUSER,
                                  SLAVE24_AWUSER,  SLAVE25_AWUSER,  SLAVE26_AWUSER,  SLAVE27_AWUSER,  SLAVE28_AWUSER,  SLAVE29_AWUSER,  SLAVE30_AWUSER,  SLAVE31_AWUSER;

  output wire                     SLAVE0_AWVALID,   SLAVE1_AWVALID,   SLAVE2_AWVALID,   SLAVE3_AWVALID,   SLAVE4_AWVALID,  SLAVE5_AWVALID,   SLAVE6_AWVALID,   SLAVE7_AWVALID,
                                  SLAVE8_AWVALID,   SLAVE9_AWVALID,   SLAVE10_AWVALID,  SLAVE11_AWVALID,  SLAVE12_AWVALID, SLAVE13_AWVALID,  SLAVE14_AWVALID,  SLAVE15_AWVALID,  
                                  SLAVE16_AWVALID,  SLAVE17_AWVALID,  SLAVE18_AWVALID,  SLAVE19_AWVALID,  SLAVE20_AWVALID, SLAVE21_AWVALID,  SLAVE22_AWVALID,   SLAVE23_AWVALID,  
                                  SLAVE24_AWVALID,  SLAVE25_AWVALID,  SLAVE26_AWVALID,  SLAVE27_AWVALID,  SLAVE28_AWVALID,  SLAVE29_AWVALID, SLAVE30_AWVALID,  SLAVE31_AWVALID;

  input  wire                     SLAVE0_AWREADY,   SLAVE1_AWREADY,   SLAVE2_AWREADY,   SLAVE3_AWREADY,   SLAVE4_AWREADY,    SLAVE5_AWREADY,   SLAVE6_AWREADY,   SLAVE7_AWREADY,
                                  SLAVE8_AWREADY,   SLAVE9_AWREADY,   SLAVE10_AWREADY,  SLAVE11_AWREADY,  SLAVE12_AWREADY,   SLAVE13_AWREADY,  SLAVE14_AWREADY,  SLAVE15_AWREADY,  
                                  SLAVE16_AWREADY,  SLAVE17_AWREADY,  SLAVE18_AWREADY,  SLAVE19_AWREADY,  SLAVE20_AWREADY,  SLAVE21_AWREADY,   SLAVE22_AWREADY,  SLAVE23_AWREADY,
                                  SLAVE24_AWREADY,  SLAVE25_AWREADY,  SLAVE26_AWREADY,  SLAVE27_AWREADY,  SLAVE28_AWREADY,  SLAVE29_AWREADY,   SLAVE30_AWREADY,  SLAVE31_AWREADY;
   
  // Slave Write Data Ports
  output wire [(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]  SLAVE0_WID,  SLAVE1_WID,  SLAVE2_WID,  SLAVE3_WID,  SLAVE4_WID,  SLAVE5_WID,  SLAVE6_WID,  SLAVE7_WID, 
                                                  SLAVE8_WID,  SLAVE9_WID,  SLAVE10_WID, SLAVE11_WID, SLAVE12_WID, SLAVE13_WID, SLAVE14_WID, SLAVE15_WID,
                                                  SLAVE16_WID, SLAVE17_WID, SLAVE18_WID, SLAVE19_WID, SLAVE20_WID, SLAVE21_WID, SLAVE22_WID, SLAVE23_WID, 
                                                  SLAVE24_WID, SLAVE25_WID, SLAVE26_WID, SLAVE27_WID, SLAVE28_WID, SLAVE29_WID, SLAVE30_WID, SLAVE31_WID;

  output wire [SLAVE0_DATA_WIDTH-1:0]      SLAVE0_WDATA;  
  output wire [SLAVE1_DATA_WIDTH-1:0]      SLAVE1_WDATA;  
  output wire [SLAVE2_DATA_WIDTH-1:0]      SLAVE2_WDATA;  
  output wire [SLAVE3_DATA_WIDTH-1:0]      SLAVE3_WDATA;  
  output wire [SLAVE4_DATA_WIDTH-1:0]      SLAVE4_WDATA;  
  output wire [SLAVE5_DATA_WIDTH-1:0]      SLAVE5_WDATA;  
  output wire [SLAVE6_DATA_WIDTH-1:0]      SLAVE6_WDATA;   
  output wire [SLAVE7_DATA_WIDTH-1:0]      SLAVE7_WDATA;  
  output wire [SLAVE8_DATA_WIDTH-1:0]      SLAVE8_WDATA;  
  output wire [SLAVE9_DATA_WIDTH-1:0]      SLAVE9_WDATA;  
  output wire [SLAVE10_DATA_WIDTH-1:0]     SLAVE10_WDATA;  
  output wire [SLAVE11_DATA_WIDTH-1:0]     SLAVE11_WDATA;  
  output wire [SLAVE12_DATA_WIDTH-1:0]     SLAVE12_WDATA;  
  output wire [SLAVE13_DATA_WIDTH-1:0]     SLAVE13_WDATA;  
  output wire [SLAVE14_DATA_WIDTH-1:0]     SLAVE14_WDATA;   
  output wire [SLAVE15_DATA_WIDTH-1:0]     SLAVE15_WDATA;  
  output wire [SLAVE16_DATA_WIDTH-1:0]     SLAVE16_WDATA;  
  output wire [SLAVE17_DATA_WIDTH-1:0]     SLAVE17_WDATA;  
  output wire [SLAVE18_DATA_WIDTH-1:0]     SLAVE18_WDATA;  
  output wire [SLAVE19_DATA_WIDTH-1:0]     SLAVE19_WDATA;  
  output wire [SLAVE20_DATA_WIDTH-1:0]     SLAVE20_WDATA;  
  output wire [SLAVE21_DATA_WIDTH-1:0]     SLAVE21_WDATA;  
  output wire [SLAVE22_DATA_WIDTH-1:0]     SLAVE22_WDATA;   
  output wire [SLAVE23_DATA_WIDTH-1:0]     SLAVE23_WDATA;  
  output wire [SLAVE24_DATA_WIDTH-1:0]     SLAVE24_WDATA;  
  output wire [SLAVE25_DATA_WIDTH-1:0]     SLAVE25_WDATA;  
  output wire [SLAVE26_DATA_WIDTH-1:0]     SLAVE26_WDATA;  
  output wire [SLAVE27_DATA_WIDTH-1:0]     SLAVE27_WDATA;  
  output wire [SLAVE28_DATA_WIDTH-1:0]     SLAVE28_WDATA;  
  output wire [SLAVE29_DATA_WIDTH-1:0]     SLAVE29_WDATA;  
  output wire [SLAVE30_DATA_WIDTH-1:0]     SLAVE30_WDATA;   
  output wire [SLAVE31_DATA_WIDTH-1:0]     SLAVE31_WDATA;
  
  
  output wire [(SLAVE0_DATA_WIDTH/8)-1:0]     SLAVE0_WSTRB;
  output wire [(SLAVE1_DATA_WIDTH/8)-1:0]     SLAVE1_WSTRB;  
  output wire [(SLAVE2_DATA_WIDTH/8)-1:0]     SLAVE2_WSTRB;  
  output wire [(SLAVE3_DATA_WIDTH/8)-1:0]     SLAVE3_WSTRB;  
  output wire [(SLAVE4_DATA_WIDTH/8)-1:0]     SLAVE4_WSTRB;  
  output wire [(SLAVE5_DATA_WIDTH/8)-1:0]     SLAVE5_WSTRB;  
  output wire [(SLAVE6_DATA_WIDTH/8)-1:0]     SLAVE6_WSTRB;  
  output wire [(SLAVE7_DATA_WIDTH/8)-1:0]     SLAVE7_WSTRB;
  output wire [(SLAVE8_DATA_WIDTH/8)-1:0]     SLAVE8_WSTRB;
  output wire [(SLAVE9_DATA_WIDTH/8)-1:0]     SLAVE9_WSTRB;  
  output wire [(SLAVE10_DATA_WIDTH/8)-1:0]    SLAVE10_WSTRB;  
  output wire [(SLAVE11_DATA_WIDTH/8)-1:0]    SLAVE11_WSTRB;  
  output wire [(SLAVE12_DATA_WIDTH/8)-1:0]    SLAVE12_WSTRB;  
  output wire [(SLAVE13_DATA_WIDTH/8)-1:0]    SLAVE13_WSTRB;  
  output wire [(SLAVE14_DATA_WIDTH/8)-1:0]    SLAVE14_WSTRB;  
  output wire [(SLAVE15_DATA_WIDTH/8)-1:0]    SLAVE15_WSTRB;
  output wire [(SLAVE16_DATA_WIDTH/8)-1:0]    SLAVE16_WSTRB;
  output wire [(SLAVE17_DATA_WIDTH/8)-1:0]    SLAVE17_WSTRB;  
  output wire [(SLAVE18_DATA_WIDTH/8)-1:0]    SLAVE18_WSTRB;  
  output wire [(SLAVE19_DATA_WIDTH/8)-1:0]    SLAVE19_WSTRB;  
  output wire [(SLAVE20_DATA_WIDTH/8)-1:0]    SLAVE20_WSTRB;  
  output wire [(SLAVE21_DATA_WIDTH/8)-1:0]    SLAVE21_WSTRB;  
  output wire [(SLAVE22_DATA_WIDTH/8)-1:0]    SLAVE22_WSTRB;  
  output wire [(SLAVE23_DATA_WIDTH/8)-1:0]    SLAVE23_WSTRB;
  output wire [(SLAVE24_DATA_WIDTH/8)-1:0]    SLAVE24_WSTRB;
  output wire [(SLAVE25_DATA_WIDTH/8)-1:0]    SLAVE25_WSTRB;  
  output wire [(SLAVE26_DATA_WIDTH/8)-1:0]    SLAVE26_WSTRB;  
  output wire [(SLAVE27_DATA_WIDTH/8)-1:0]    SLAVE27_WSTRB;  
  output wire [(SLAVE28_DATA_WIDTH/8)-1:0]    SLAVE28_WSTRB;  
  output wire [(SLAVE29_DATA_WIDTH/8)-1:0]    SLAVE29_WSTRB;  
  output wire [(SLAVE30_DATA_WIDTH/8)-1:0]    SLAVE30_WSTRB;  
  output wire [(SLAVE31_DATA_WIDTH/8)-1:0]    SLAVE31_WSTRB;
  
  
  output wire                         SLAVE0_WLAST,  SLAVE1_WLAST,  SLAVE2_WLAST,  SLAVE3_WLAST,  SLAVE4_WLAST,  SLAVE5_WLAST,  SLAVE6_WLAST,  SLAVE7_WLAST, 
                                      SLAVE8_WLAST,  SLAVE9_WLAST,  SLAVE10_WLAST, SLAVE11_WLAST, SLAVE12_WLAST, SLAVE13_WLAST, SLAVE14_WLAST, SLAVE15_WLAST, 
                                      SLAVE16_WLAST, SLAVE17_WLAST, SLAVE18_WLAST, SLAVE19_WLAST, SLAVE20_WLAST, SLAVE21_WLAST, SLAVE22_WLAST, SLAVE23_WLAST, 
                                      SLAVE24_WLAST, SLAVE25_WLAST, SLAVE26_WLAST, SLAVE27_WLAST, SLAVE28_WLAST, SLAVE29_WLAST, SLAVE30_WLAST, SLAVE31_WLAST;
                                      
  output wire [USER_WIDTH-1:0]        SLAVE0_WUSER,  SLAVE1_WUSER,  SLAVE2_WUSER,  SLAVE3_WUSER,  SLAVE4_WUSER,  SLAVE5_WUSER,  SLAVE6_WUSER,  SLAVE7_WUSER, 
                                      SLAVE8_WUSER,  SLAVE9_WUSER,  SLAVE10_WUSER, SLAVE11_WUSER, SLAVE12_WUSER, SLAVE13_WUSER, SLAVE14_WUSER, SLAVE15_WUSER, 
                                      SLAVE16_WUSER, SLAVE17_WUSER, SLAVE18_WUSER, SLAVE19_WUSER, SLAVE20_WUSER, SLAVE21_WUSER, SLAVE22_WUSER, SLAVE23_WUSER, 
                                      SLAVE24_WUSER, SLAVE25_WUSER, SLAVE26_WUSER, SLAVE27_WUSER, SLAVE28_WUSER, SLAVE29_WUSER, SLAVE30_WUSER, SLAVE31_WUSER;
                                      
  output wire                         SLAVE0_WVALID,  SLAVE1_WVALID,  SLAVE2_WVALID,  SLAVE3_WVALID,  SLAVE4_WVALID,  SLAVE5_WVALID,  SLAVE6_WVALID,  SLAVE7_WVALID, 
                                      SLAVE8_WVALID,  SLAVE9_WVALID,  SLAVE10_WVALID, SLAVE11_WVALID, SLAVE12_WVALID, SLAVE13_WVALID, SLAVE14_WVALID, SLAVE15_WVALID, 
                                      SLAVE16_WVALID, SLAVE17_WVALID, SLAVE18_WVALID, SLAVE19_WVALID, SLAVE20_WVALID, SLAVE21_WVALID, SLAVE22_WVALID, SLAVE23_WVALID, 
                                      SLAVE24_WVALID, SLAVE25_WVALID, SLAVE26_WVALID, SLAVE27_WVALID, SLAVE28_WVALID, SLAVE29_WVALID, SLAVE30_WVALID, SLAVE31_WVALID;
                                      
  input  wire                         SLAVE0_WREADY,  SLAVE1_WREADY,  SLAVE2_WREADY,  SLAVE3_WREADY,  SLAVE4_WREADY,  SLAVE5_WREADY,  SLAVE6_WREADY,  SLAVE7_WREADY, 
                                      SLAVE8_WREADY,  SLAVE9_WREADY,  SLAVE10_WREADY, SLAVE11_WREADY, SLAVE12_WREADY, SLAVE13_WREADY, SLAVE14_WREADY, SLAVE15_WREADY, 
                                      SLAVE16_WREADY, SLAVE17_WREADY, SLAVE18_WREADY, SLAVE19_WREADY, SLAVE20_WREADY, SLAVE21_WREADY, SLAVE22_WREADY, SLAVE23_WREADY, 
                                      SLAVE24_WREADY, SLAVE25_WREADY, SLAVE26_WREADY, SLAVE27_WREADY, SLAVE28_WREADY, SLAVE29_WREADY, SLAVE30_WREADY, SLAVE31_WREADY;

  // Slave Write Response Ports
  input  wire [(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE0_BID,  SLAVE1_BID,  SLAVE2_BID,  SLAVE3_BID,  SLAVE4_BID,  SLAVE5_BID,  SLAVE6_BID,  SLAVE7_BID, 
                                                    SLAVE8_BID,  SLAVE9_BID,  SLAVE10_BID, SLAVE11_BID, SLAVE12_BID, SLAVE13_BID, SLAVE14_BID, SLAVE15_BID, 
                                                    SLAVE16_BID, SLAVE17_BID, SLAVE18_BID, SLAVE19_BID, SLAVE20_BID, SLAVE21_BID, SLAVE22_BID, SLAVE23_BID, 
                                                    SLAVE24_BID, SLAVE25_BID, SLAVE26_BID, SLAVE27_BID, SLAVE28_BID, SLAVE29_BID, SLAVE30_BID, SLAVE31_BID;
                                                    
  input  wire [1:0]                                 SLAVE0_BRESP,  SLAVE1_BRESP,  SLAVE2_BRESP,  SLAVE3_BRESP,  SLAVE4_BRESP,  SLAVE5_BRESP,  SLAVE6_BRESP,  SLAVE7_BRESP, 
                                                    SLAVE8_BRESP,  SLAVE9_BRESP,  SLAVE10_BRESP, SLAVE11_BRESP, SLAVE12_BRESP, SLAVE13_BRESP, SLAVE14_BRESP, SLAVE15_BRESP, 
                                                    SLAVE16_BRESP, SLAVE17_BRESP, SLAVE18_BRESP, SLAVE19_BRESP, SLAVE20_BRESP, SLAVE21_BRESP, SLAVE22_BRESP, SLAVE23_BRESP, 
                                                    SLAVE24_BRESP, SLAVE25_BRESP, SLAVE26_BRESP, SLAVE27_BRESP, SLAVE28_BRESP, SLAVE29_BRESP, SLAVE30_BRESP, SLAVE31_BRESP;
                            
  input  wire [USER_WIDTH-1:0]                      SLAVE0_BUSER,  SLAVE1_BUSER,  SLAVE2_BUSER,  SLAVE3_BUSER,  SLAVE4_BUSER,  SLAVE5_BUSER,  SLAVE6_BUSER,  SLAVE7_BUSER, 
                                                    SLAVE8_BUSER,  SLAVE9_BUSER,  SLAVE10_BUSER, SLAVE11_BUSER, SLAVE12_BUSER, SLAVE13_BUSER, SLAVE14_BUSER, SLAVE15_BUSER, 
                                                    SLAVE16_BUSER, SLAVE17_BUSER, SLAVE18_BUSER, SLAVE19_BUSER, SLAVE20_BUSER, SLAVE21_BUSER, SLAVE22_BUSER, SLAVE23_BUSER, 
                                                    SLAVE24_BUSER, SLAVE25_BUSER, SLAVE26_BUSER, SLAVE27_BUSER, SLAVE28_BUSER, SLAVE29_BUSER, SLAVE30_BUSER, SLAVE31_BUSER;
                                                    
  input  wire                                       SLAVE0_BVALID,  SLAVE1_BVALID,  SLAVE2_BVALID,  SLAVE3_BVALID,  SLAVE4_BVALID,  SLAVE5_BVALID,  SLAVE6_BVALID,  SLAVE7_BVALID, 
                                                    SLAVE8_BVALID,  SLAVE9_BVALID,  SLAVE10_BVALID, SLAVE11_BVALID, SLAVE12_BVALID, SLAVE13_BVALID, SLAVE14_BVALID, SLAVE15_BVALID, 
                                                    SLAVE16_BVALID, SLAVE17_BVALID, SLAVE18_BVALID, SLAVE19_BVALID, SLAVE20_BVALID, SLAVE21_BVALID, SLAVE22_BVALID, SLAVE23_BVALID, 
                                                    SLAVE24_BVALID, SLAVE25_BVALID, SLAVE26_BVALID, SLAVE27_BVALID, SLAVE28_BVALID, SLAVE29_BVALID, SLAVE30_BVALID, SLAVE31_BVALID;

  output wire                                       SLAVE0_BREADY,  SLAVE1_BREADY,  SLAVE2_BREADY,  SLAVE3_BREADY,  SLAVE4_BREADY,  SLAVE5_BREADY,  SLAVE6_BREADY,  SLAVE7_BREADY, 
                                                    SLAVE8_BREADY,  SLAVE9_BREADY,  SLAVE10_BREADY, SLAVE11_BREADY, SLAVE12_BREADY, SLAVE13_BREADY, SLAVE14_BREADY, SLAVE15_BREADY, 
                                                    SLAVE16_BREADY, SLAVE17_BREADY, SLAVE18_BREADY, SLAVE19_BREADY, SLAVE20_BREADY, SLAVE21_BREADY, SLAVE22_BREADY, SLAVE23_BREADY, 
                                                    SLAVE24_BREADY, SLAVE25_BREADY, SLAVE26_BREADY, SLAVE27_BREADY, SLAVE28_BREADY, SLAVE29_BREADY, SLAVE30_BREADY, SLAVE31_BREADY;
   
  // Slave Read Address Port
  output wire [(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE0_ARID,  SLAVE1_ARID,  SLAVE2_ARID,  SLAVE3_ARID,  SLAVE4_ARID,  SLAVE5_ARID,  SLAVE6_ARID,  SLAVE7_ARID, 
                                                    SLAVE8_ARID,  SLAVE9_ARID,  SLAVE10_ARID, SLAVE11_ARID, SLAVE12_ARID, SLAVE13_ARID, SLAVE14_ARID, SLAVE15_ARID, 
                                                    SLAVE16_ARID, SLAVE17_ARID, SLAVE18_ARID, SLAVE19_ARID, SLAVE20_ARID, SLAVE21_ARID, SLAVE22_ARID, SLAVE23_ARID, 
                                                    SLAVE24_ARID, SLAVE25_ARID, SLAVE26_ARID, SLAVE27_ARID, SLAVE28_ARID, SLAVE29_ARID, SLAVE30_ARID, SLAVE31_ARID;
  
  
  
  output wire [ADDR_WIDTH-1:0]      SLAVE0_ARADDR,  SLAVE1_ARADDR,  SLAVE2_ARADDR,  SLAVE3_ARADDR,  SLAVE4_ARADDR,  SLAVE5_ARADDR,  SLAVE6_ARADDR,  SLAVE7_ARADDR, 
                                    SLAVE8_ARADDR,  SLAVE9_ARADDR,  SLAVE10_ARADDR, SLAVE11_ARADDR, SLAVE12_ARADDR, SLAVE13_ARADDR, SLAVE14_ARADDR, SLAVE15_ARADDR, 
                                    SLAVE16_ARADDR, SLAVE17_ARADDR, SLAVE18_ARADDR, SLAVE19_ARADDR, SLAVE20_ARADDR, SLAVE21_ARADDR, SLAVE22_ARADDR, SLAVE23_ARADDR, 
                                    SLAVE24_ARADDR, SLAVE25_ARADDR, SLAVE26_ARADDR, SLAVE27_ARADDR, SLAVE28_ARADDR, SLAVE29_ARADDR, SLAVE30_ARADDR, SLAVE31_ARADDR;


  output wire [7:0]                 SLAVE0_ARLEN,  SLAVE1_ARLEN,  SLAVE2_ARLEN,  SLAVE3_ARLEN,  SLAVE4_ARLEN,  SLAVE5_ARLEN,  SLAVE6_ARLEN,  SLAVE7_ARLEN, 
                                    SLAVE8_ARLEN,  SLAVE9_ARLEN,  SLAVE10_ARLEN, SLAVE11_ARLEN, SLAVE12_ARLEN, SLAVE13_ARLEN, SLAVE14_ARLEN, SLAVE15_ARLEN, 
                                    SLAVE16_ARLEN, SLAVE17_ARLEN, SLAVE18_ARLEN, SLAVE19_ARLEN, SLAVE20_ARLEN, SLAVE21_ARLEN, SLAVE22_ARLEN, SLAVE23_ARLEN, 
                                    SLAVE24_ARLEN, SLAVE25_ARLEN, SLAVE26_ARLEN, SLAVE27_ARLEN, SLAVE28_ARLEN, SLAVE29_ARLEN, SLAVE30_ARLEN, SLAVE31_ARLEN;


  output wire [2:0]                 SLAVE0_ARSIZE,  SLAVE1_ARSIZE,  SLAVE2_ARSIZE,  SLAVE3_ARSIZE,  SLAVE4_ARSIZE,  SLAVE5_ARSIZE,  SLAVE6_ARSIZE,  SLAVE7_ARSIZE, 
                                    SLAVE8_ARSIZE,  SLAVE9_ARSIZE,  SLAVE10_ARSIZE, SLAVE11_ARSIZE, SLAVE12_ARSIZE, SLAVE13_ARSIZE, SLAVE14_ARSIZE, SLAVE15_ARSIZE, 
                                    SLAVE16_ARSIZE, SLAVE17_ARSIZE, SLAVE18_ARSIZE, SLAVE19_ARSIZE, SLAVE20_ARSIZE, SLAVE21_ARSIZE, SLAVE22_ARSIZE, SLAVE23_ARSIZE, 
                                    SLAVE24_ARSIZE, SLAVE25_ARSIZE, SLAVE26_ARSIZE, SLAVE27_ARSIZE, SLAVE28_ARSIZE, SLAVE29_ARSIZE, SLAVE30_ARSIZE, SLAVE31_ARSIZE;


  output wire [1:0]                 SLAVE0_ARBURST,  SLAVE1_ARBURST,  SLAVE2_ARBURST,  SLAVE3_ARBURST,  SLAVE4_ARBURST,  SLAVE5_ARBURST,  SLAVE6_ARBURST,  SLAVE7_ARBURST, 
                                    SLAVE8_ARBURST,  SLAVE9_ARBURST,  SLAVE10_ARBURST, SLAVE11_ARBURST, SLAVE12_ARBURST, SLAVE13_ARBURST, SLAVE14_ARBURST, SLAVE15_ARBURST, 
                                    SLAVE16_ARBURST, SLAVE17_ARBURST, SLAVE18_ARBURST, SLAVE19_ARBURST, SLAVE20_ARBURST, SLAVE21_ARBURST, SLAVE22_ARBURST, SLAVE23_ARBURST, 
                                    SLAVE24_ARBURST, SLAVE25_ARBURST, SLAVE26_ARBURST, SLAVE27_ARBURST, SLAVE28_ARBURST, SLAVE29_ARBURST, SLAVE30_ARBURST, SLAVE31_ARBURST;


  output wire [1:0]                 SLAVE0_ARLOCK,  SLAVE1_ARLOCK,  SLAVE2_ARLOCK,  SLAVE3_ARLOCK,  SLAVE4_ARLOCK,  SLAVE5_ARLOCK,  SLAVE6_ARLOCK,  SLAVE7_ARLOCK, 
                                    SLAVE8_ARLOCK,  SLAVE9_ARLOCK,  SLAVE10_ARLOCK, SLAVE11_ARLOCK, SLAVE12_ARLOCK, SLAVE13_ARLOCK, SLAVE14_ARLOCK, SLAVE15_ARLOCK, 
                                    SLAVE16_ARLOCK, SLAVE17_ARLOCK, SLAVE18_ARLOCK, SLAVE19_ARLOCK, SLAVE20_ARLOCK, SLAVE21_ARLOCK, SLAVE22_ARLOCK, SLAVE23_ARLOCK, 
                                    SLAVE24_ARLOCK, SLAVE25_ARLOCK, SLAVE26_ARLOCK, SLAVE27_ARLOCK, SLAVE28_ARLOCK, SLAVE29_ARLOCK, SLAVE30_ARLOCK, SLAVE31_ARLOCK;


  output wire [3:0]                 SLAVE0_ARCACHE,  SLAVE1_ARCACHE,  SLAVE2_ARCACHE,  SLAVE3_ARCACHE,  SLAVE4_ARCACHE,  SLAVE5_ARCACHE,  SLAVE6_ARCACHE,  SLAVE7_ARCACHE, 
                                    SLAVE8_ARCACHE,  SLAVE9_ARCACHE,  SLAVE10_ARCACHE, SLAVE11_ARCACHE, SLAVE12_ARCACHE, SLAVE13_ARCACHE, SLAVE14_ARCACHE, SLAVE15_ARCACHE, 
                                    SLAVE16_ARCACHE, SLAVE17_ARCACHE, SLAVE18_ARCACHE, SLAVE19_ARCACHE, SLAVE20_ARCACHE, SLAVE21_ARCACHE, SLAVE22_ARCACHE, SLAVE23_ARCACHE, 
                                    SLAVE24_ARCACHE, SLAVE25_ARCACHE, SLAVE26_ARCACHE, SLAVE27_ARCACHE, SLAVE28_ARCACHE, SLAVE29_ARCACHE, SLAVE30_ARCACHE, SLAVE31_ARCACHE;


  output wire [2:0]                 SLAVE0_ARPROT,  SLAVE1_ARPROT,  SLAVE2_ARPROT,  SLAVE3_ARPROT,  SLAVE4_ARPROT,  SLAVE5_ARPROT,  SLAVE6_ARPROT,  SLAVE7_ARPROT, 
                                    SLAVE8_ARPROT,  SLAVE9_ARPROT,  SLAVE10_ARPROT, SLAVE11_ARPROT, SLAVE12_ARPROT, SLAVE13_ARPROT, SLAVE14_ARPROT, SLAVE15_ARPROT, 
                                    SLAVE16_ARPROT, SLAVE17_ARPROT, SLAVE18_ARPROT, SLAVE19_ARPROT, SLAVE20_ARPROT, SLAVE21_ARPROT, SLAVE22_ARPROT, SLAVE23_ARPROT, 
                                    SLAVE24_ARPROT, SLAVE25_ARPROT, SLAVE26_ARPROT, SLAVE27_ARPROT, SLAVE28_ARPROT, SLAVE29_ARPROT, SLAVE30_ARPROT, SLAVE31_ARPROT;


  output wire [3:0]                 SLAVE0_ARREGION,  SLAVE1_ARREGION,  SLAVE2_ARREGION,  SLAVE3_ARREGION,  SLAVE4_ARREGION,  SLAVE5_ARREGION,  SLAVE6_ARREGION,  SLAVE7_ARREGION, 
                                    SLAVE8_ARREGION,  SLAVE9_ARREGION,  SLAVE10_ARREGION, SLAVE11_ARREGION, SLAVE12_ARREGION, SLAVE13_ARREGION, SLAVE14_ARREGION, SLAVE15_ARREGION, 
                                    SLAVE16_ARREGION, SLAVE17_ARREGION, SLAVE18_ARREGION, SLAVE19_ARREGION, SLAVE20_ARREGION, SLAVE21_ARREGION, SLAVE22_ARREGION, SLAVE23_ARREGION, 
                                    SLAVE24_ARREGION, SLAVE25_ARREGION, SLAVE26_ARREGION, SLAVE27_ARREGION, SLAVE28_ARREGION, SLAVE29_ARREGION, SLAVE30_ARREGION, SLAVE31_ARREGION;


  output wire [3:0]                 SLAVE0_ARQOS,  SLAVE1_ARQOS,  SLAVE2_ARQOS,  SLAVE3_ARQOS,  SLAVE4_ARQOS,  SLAVE5_ARQOS,  SLAVE6_ARQOS,  SLAVE7_ARQOS, 
                                    SLAVE8_ARQOS,  SLAVE9_ARQOS,  SLAVE10_ARQOS, SLAVE11_ARQOS, SLAVE12_ARQOS, SLAVE13_ARQOS, SLAVE14_ARQOS, SLAVE15_ARQOS, 
                                    SLAVE16_ARQOS, SLAVE17_ARQOS, SLAVE18_ARQOS, SLAVE19_ARQOS, SLAVE20_ARQOS, SLAVE21_ARQOS, SLAVE22_ARQOS, SLAVE23_ARQOS, 
                                    SLAVE24_ARQOS, SLAVE25_ARQOS, SLAVE26_ARQOS, SLAVE27_ARQOS, SLAVE28_ARQOS, SLAVE29_ARQOS, SLAVE30_ARQOS, SLAVE31_ARQOS;

  output wire [USER_WIDTH-1:0]      SLAVE0_ARUSER,  SLAVE1_ARUSER,  SLAVE2_ARUSER,  SLAVE3_ARUSER,  SLAVE4_ARUSER,  SLAVE5_ARUSER,  SLAVE6_ARUSER,  SLAVE7_ARUSER, 
                                    SLAVE8_ARUSER,  SLAVE9_ARUSER,  SLAVE10_ARUSER, SLAVE11_ARUSER, SLAVE12_ARUSER, SLAVE13_ARUSER, SLAVE14_ARUSER, SLAVE15_ARUSER, 
                                    SLAVE16_ARUSER, SLAVE17_ARUSER, SLAVE18_ARUSER, SLAVE19_ARUSER, SLAVE20_ARUSER, SLAVE21_ARUSER, SLAVE22_ARUSER, SLAVE23_ARUSER, 
                                    SLAVE24_ARUSER, SLAVE25_ARUSER, SLAVE26_ARUSER, SLAVE27_ARUSER, SLAVE28_ARUSER, SLAVE29_ARUSER, SLAVE30_ARUSER, SLAVE31_ARUSER;


  output wire                       SLAVE0_ARVALID,  SLAVE1_ARVALID,  SLAVE2_ARVALID,  SLAVE3_ARVALID,  SLAVE4_ARVALID,  SLAVE5_ARVALID,  SLAVE6_ARVALID,  SLAVE7_ARVALID, 
                                    SLAVE8_ARVALID,  SLAVE9_ARVALID,  SLAVE10_ARVALID, SLAVE11_ARVALID, SLAVE12_ARVALID, SLAVE13_ARVALID, SLAVE14_ARVALID, SLAVE15_ARVALID, 
                                    SLAVE16_ARVALID, SLAVE17_ARVALID, SLAVE18_ARVALID, SLAVE19_ARVALID, SLAVE20_ARVALID, SLAVE21_ARVALID, SLAVE22_ARVALID, SLAVE23_ARVALID, 
                                    SLAVE24_ARVALID, SLAVE25_ARVALID, SLAVE26_ARVALID, SLAVE27_ARVALID, SLAVE28_ARVALID, SLAVE29_ARVALID, SLAVE30_ARVALID, SLAVE31_ARVALID;

  
  input  wire                       SLAVE0_ARREADY,  SLAVE1_ARREADY,  SLAVE2_ARREADY,  SLAVE3_ARREADY,  SLAVE4_ARREADY,  SLAVE5_ARREADY,  SLAVE6_ARREADY,  SLAVE7_ARREADY, 
                                    SLAVE8_ARREADY,  SLAVE9_ARREADY,  SLAVE10_ARREADY, SLAVE11_ARREADY, SLAVE12_ARREADY, SLAVE13_ARREADY, SLAVE14_ARREADY, SLAVE15_ARREADY, 
                                    SLAVE16_ARREADY, SLAVE17_ARREADY, SLAVE18_ARREADY, SLAVE19_ARREADY, SLAVE20_ARREADY, SLAVE21_ARREADY, SLAVE22_ARREADY, SLAVE23_ARREADY, 
                                    SLAVE24_ARREADY, SLAVE25_ARREADY, SLAVE26_ARREADY, SLAVE27_ARREADY, SLAVE28_ARREADY, SLAVE29_ARREADY, SLAVE30_ARREADY, SLAVE31_ARREADY;


  // Slave Read Data Ports
  input  wire [(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE0_RID,  SLAVE1_RID,  SLAVE2_RID,  SLAVE3_RID,  SLAVE4_RID,  SLAVE5_RID,  SLAVE6_RID,  SLAVE7_RID, 
                                                    SLAVE8_RID,  SLAVE9_RID,  SLAVE10_RID, SLAVE11_RID, SLAVE12_RID, SLAVE13_RID, SLAVE14_RID, SLAVE15_RID, 
                                                    SLAVE16_RID, SLAVE17_RID, SLAVE18_RID, SLAVE19_RID, SLAVE20_RID, SLAVE21_RID, SLAVE22_RID, SLAVE23_RID, 
                                                    SLAVE24_RID, SLAVE25_RID, SLAVE26_RID, SLAVE27_RID, SLAVE28_RID, SLAVE29_RID, SLAVE30_RID, SLAVE31_RID;
                                                    
  input  wire [SLAVE0_DATA_WIDTH-1:0]    SLAVE0_RDATA;
  input  wire [SLAVE1_DATA_WIDTH-1:0]    SLAVE1_RDATA;
  input  wire [SLAVE2_DATA_WIDTH-1:0]    SLAVE2_RDATA;
  input  wire [SLAVE3_DATA_WIDTH-1:0]    SLAVE3_RDATA;
  input  wire [SLAVE4_DATA_WIDTH-1:0]    SLAVE4_RDATA;
  input  wire [SLAVE5_DATA_WIDTH-1:0]    SLAVE5_RDATA;
  input  wire [SLAVE6_DATA_WIDTH-1:0]    SLAVE6_RDATA;
  input  wire [SLAVE7_DATA_WIDTH-1:0]    SLAVE7_RDATA;
  input  wire [SLAVE8_DATA_WIDTH-1:0]    SLAVE8_RDATA;
  input  wire [SLAVE9_DATA_WIDTH-1:0]    SLAVE9_RDATA;
  input  wire [SLAVE10_DATA_WIDTH-1:0]   SLAVE10_RDATA;
  input  wire [SLAVE11_DATA_WIDTH-1:0]   SLAVE11_RDATA;
  input  wire [SLAVE12_DATA_WIDTH-1:0]   SLAVE12_RDATA;
  input  wire [SLAVE13_DATA_WIDTH-1:0]   SLAVE13_RDATA;
  input  wire [SLAVE14_DATA_WIDTH-1:0]   SLAVE14_RDATA;
  input  wire [SLAVE15_DATA_WIDTH-1:0]   SLAVE15_RDATA;
  input  wire [SLAVE16_DATA_WIDTH-1:0]   SLAVE16_RDATA;
  input  wire [SLAVE17_DATA_WIDTH-1:0]   SLAVE17_RDATA;
  input  wire [SLAVE18_DATA_WIDTH-1:0]   SLAVE18_RDATA;
  input  wire [SLAVE19_DATA_WIDTH-1:0]   SLAVE19_RDATA;
  input  wire [SLAVE20_DATA_WIDTH-1:0]   SLAVE20_RDATA;
  input  wire [SLAVE21_DATA_WIDTH-1:0]   SLAVE21_RDATA;
  input  wire [SLAVE22_DATA_WIDTH-1:0]   SLAVE22_RDATA;
  input  wire [SLAVE23_DATA_WIDTH-1:0]   SLAVE23_RDATA;
  input  wire [SLAVE24_DATA_WIDTH-1:0]   SLAVE24_RDATA;
  input  wire [SLAVE25_DATA_WIDTH-1:0]   SLAVE25_RDATA;
  input  wire [SLAVE26_DATA_WIDTH-1:0]   SLAVE26_RDATA;
  input  wire [SLAVE27_DATA_WIDTH-1:0]   SLAVE27_RDATA;
  input  wire [SLAVE28_DATA_WIDTH-1:0]   SLAVE28_RDATA;
  input  wire [SLAVE29_DATA_WIDTH-1:0]   SLAVE29_RDATA;
  input  wire [SLAVE30_DATA_WIDTH-1:0]   SLAVE30_RDATA;
  input  wire [SLAVE31_DATA_WIDTH-1:0]   SLAVE31_RDATA;
  
  
  input  wire [1:0]                 SLAVE0_RRESP,  SLAVE1_RRESP,  SLAVE2_RRESP,  SLAVE3_RRESP,  SLAVE4_RRESP,  SLAVE5_RRESP,  SLAVE6_RRESP,  SLAVE7_RRESP,
                                    SLAVE8_RRESP,  SLAVE9_RRESP,  SLAVE10_RRESP, SLAVE11_RRESP, SLAVE12_RRESP, SLAVE13_RRESP, SLAVE14_RRESP, SLAVE15_RRESP, 
                                    SLAVE16_RRESP, SLAVE17_RRESP, SLAVE18_RRESP, SLAVE19_RRESP, SLAVE20_RRESP, SLAVE21_RRESP, SLAVE22_RRESP, SLAVE23_RRESP, 
                                    SLAVE24_RRESP, SLAVE25_RRESP, SLAVE26_RRESP, SLAVE27_RRESP, SLAVE28_RRESP, SLAVE29_RRESP, SLAVE30_RRESP, SLAVE31_RRESP;

  input  wire                       SLAVE0_RLAST,  SLAVE1_RLAST,  SLAVE2_RLAST,  SLAVE3_RLAST,  SLAVE4_RLAST,  SLAVE5_RLAST,  SLAVE6_RLAST,  SLAVE7_RLAST,
                                    SLAVE8_RLAST,  SLAVE9_RLAST,  SLAVE10_RLAST, SLAVE11_RLAST, SLAVE12_RLAST, SLAVE13_RLAST, SLAVE14_RLAST, SLAVE15_RLAST, 
                                    SLAVE16_RLAST, SLAVE17_RLAST, SLAVE18_RLAST, SLAVE19_RLAST, SLAVE20_RLAST, SLAVE21_RLAST, SLAVE22_RLAST, SLAVE23_RLAST, 
                                    SLAVE24_RLAST, SLAVE25_RLAST, SLAVE26_RLAST, SLAVE27_RLAST, SLAVE28_RLAST, SLAVE29_RLAST, SLAVE30_RLAST, SLAVE31_RLAST;
                                                    
                                                    
  input  wire [USER_WIDTH-1:0]      SLAVE0_RUSER,  SLAVE1_RUSER,  SLAVE2_RUSER,  SLAVE3_RUSER,  SLAVE4_RUSER,  SLAVE5_RUSER,  SLAVE6_RUSER,  SLAVE7_RUSER,
                                    SLAVE8_RUSER,  SLAVE9_RUSER,  SLAVE10_RUSER, SLAVE11_RUSER, SLAVE12_RUSER, SLAVE13_RUSER, SLAVE14_RUSER, SLAVE15_RUSER, 
                                    SLAVE16_RUSER, SLAVE17_RUSER, SLAVE18_RUSER, SLAVE19_RUSER, SLAVE20_RUSER, SLAVE21_RUSER, SLAVE22_RUSER, SLAVE23_RUSER, 
                                    SLAVE24_RUSER, SLAVE25_RUSER, SLAVE26_RUSER, SLAVE27_RUSER, SLAVE28_RUSER, SLAVE29_RUSER, SLAVE30_RUSER, SLAVE31_RUSER;
                                                    
                                                    
  input  wire                       SLAVE0_RVALID,  SLAVE1_RVALID,  SLAVE2_RVALID,  SLAVE3_RVALID,  SLAVE4_RVALID,  SLAVE5_RVALID,  SLAVE6_RVALID,   SLAVE7_RVALID,
                                    SLAVE8_RVALID,  SLAVE9_RVALID,  SLAVE10_RVALID, SLAVE11_RVALID, SLAVE12_RVALID, SLAVE13_RVALID, SLAVE14_RVALID, SLAVE15_RVALID, 
                                    SLAVE16_RVALID, SLAVE17_RVALID, SLAVE18_RVALID, SLAVE19_RVALID, SLAVE20_RVALID, SLAVE21_RVALID, SLAVE22_RVALID, SLAVE23_RVALID, 
                                    SLAVE24_RVALID, SLAVE25_RVALID, SLAVE26_RVALID, SLAVE27_RVALID, SLAVE28_RVALID, SLAVE29_RVALID, SLAVE30_RVALID, SLAVE31_RVALID;
                                                    
                                                    
  output wire                       SLAVE0_RREADY,  SLAVE1_RREADY,  SLAVE2_RREADY,  SLAVE3_RREADY,  SLAVE4_RREADY,  SLAVE5_RREADY,  SLAVE6_RREADY,  SLAVE7_RREADY,
                                    SLAVE8_RREADY,  SLAVE9_RREADY,  SLAVE10_RREADY, SLAVE11_RREADY, SLAVE12_RREADY, SLAVE13_RREADY, SLAVE14_RREADY, SLAVE15_RREADY, 
                                    SLAVE16_RREADY, SLAVE17_RREADY, SLAVE18_RREADY, SLAVE19_RREADY, SLAVE20_RREADY, SLAVE21_RREADY, SLAVE22_RREADY, SLAVE23_RREADY, 
                                    SLAVE24_RREADY, SLAVE25_RREADY, SLAVE26_RREADY, SLAVE27_RREADY, SLAVE28_RREADY, SLAVE29_RREADY, SLAVE30_RREADY, SLAVE31_RREADY;
   
  //==================================================================================================================================
  // Variable Declarations
  //==================================================================================================================================  

  //====================== Slave Read Address Ports  ================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0] slaveARID;
  wire [NUM_SLAVES*ADDR_WIDTH-1:0]                   slaveARADDR;
  wire [NUM_SLAVES*8-1:0]                            slaveARLEN;
  wire [NUM_SLAVES*3-1:0]                            slaveARSIZE;
  wire [NUM_SLAVES*2-1:0]                            slaveARBURST;
  wire [NUM_SLAVES*2-1:0]                            slaveARLOCK;
  wire [NUM_SLAVES*4-1:0]                            slaveARCACHE;
  wire [NUM_SLAVES*3-1:0]                            slaveARPROT;
  wire [NUM_SLAVES*4-1:0]                            slaveARREGION;
  wire [NUM_SLAVES*4-1:0]                            slaveARQOS;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                   slaveARUSER;
  wire [NUM_SLAVES-1:0]                              slaveARVALID;
  wire [NUM_SLAVES-1:0]                              slaveARREADY;

  //====================== Slave Read Data Ports  ====================================================//
  wire [NUM_SLAVES-1:0]                               slaveRVALID;
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]  slaveRID;
  wire [NUM_SLAVES*DATA_WIDTH-1:0]                    slaveRDATA;
  wire [NUM_SLAVES*2-1:0]                             slaveRRESP;
  wire [NUM_SLAVES-1:0]                               slaveRLAST;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                    slaveRUSER;
    
  wire [NUM_SLAVES-1:0]                               slaveRREADY;

  //====================== Slave Write Address Ports  ====================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]  slaveAWID;
  wire [NUM_SLAVES*ADDR_WIDTH-1:0]                    slaveAWADDR;
  wire [NUM_SLAVES*8-1:0]                             slaveAWLEN;
  wire [NUM_SLAVES*3-1:0]                             slaveAWSIZE;
  wire [NUM_SLAVES*2-1:0]                             slaveAWBURST;
  wire [NUM_SLAVES*2-1:0]                             slaveAWLOCK;
  wire [NUM_SLAVES*4-1:0]                             slaveAWCACHE;
  wire [NUM_SLAVES*3-1:0]                             slaveAWPROT;
  wire [NUM_SLAVES*4-1:0]                             slaveAWREGION;
  wire [NUM_SLAVES*4-1:0]                             slaveAWQOS;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                    slaveAWUSER;
  wire [NUM_SLAVES-1:0]                               slaveAWVALID;
  wire [NUM_SLAVES-1:0]                               slaveAWREADY;

  //====================== Slave Write Data Ports  ====================================================//
  wire [NUM_SLAVES*DATA_WIDTH-1:0]                    slaveWDATA;
  wire [NUM_SLAVES*DATA_WIDTH/8-1:0]                  slaveWSTRB;
  wire [NUM_SLAVES-1:0]                               slaveWLAST;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                    slaveWUSER;
  wire [NUM_SLAVES-1:0]                               slaveWVALID;
  wire [NUM_SLAVES-1:0]                               slaveWREADY;

  //====================== Slave Write Response Ports  ====================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]  slaveBID;
  wire [NUM_SLAVES*2-1:0]                             slaveBRESP;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                    slaveBUSER;
  wire [NUM_SLAVES-1:0]                               slaveBVALID;
  wire [NUM_SLAVES-1:0]                               slaveBREADY;


  //====================== Slave Read Address Ports  ================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE_ARID;
  wire [NUM_SLAVES*ADDR_WIDTH-1:0]                      SLAVE_ARADDR;
  wire [NUM_SLAVES*8-1:0]                               SLAVE_ARLEN;
  wire [NUM_SLAVES*3-1:0]                               SLAVE_ARSIZE;
  wire [NUM_SLAVES*2-1:0]                               SLAVE_ARBURST;
  wire [NUM_SLAVES*2-1:0]                               SLAVE_ARLOCK;
  wire [NUM_SLAVES*4-1:0]                               SLAVE_ARCACHE;
  wire [NUM_SLAVES*3-1:0]                               SLAVE_ARPROT;
  wire [NUM_SLAVES*4-1:0]                               SLAVE_ARREGION;
  wire [NUM_SLAVES*4-1:0]                               SLAVE_ARQOS;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                      SLAVE_ARUSER;
  wire [NUM_SLAVES-1:0]                                 SLAVE_ARVALID;
  wire [NUM_SLAVES-1:0]                                 SLAVE_ARREADY;

  //====================== Slave Read Data Ports  ====================================================//
  wire [NUM_SLAVES-1:0]                                 SLAVE_RVALID;
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE_RID;
  wire [SLAVE_DATA_WIDTH_PORT-1:0]                      SLAVE_RDATA;
  wire [NUM_SLAVES*2-1:0]                               SLAVE_RRESP;
  wire [NUM_SLAVES-1:0]                                 SLAVE_RLAST;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                      SLAVE_RUSER;    
  wire [NUM_SLAVES-1:0]                                 SLAVE_RREADY;

  //====================== Slave Write Address Ports  ====================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE_AWID;
  wire [NUM_SLAVES*ADDR_WIDTH-1:0]                      SLAVE_AWADDR;
  wire [NUM_SLAVES*8-1:0]                               SLAVE_AWLEN;
  wire [NUM_SLAVES*3-1:0]                               SLAVE_AWSIZE;
  wire [NUM_SLAVES*2-1:0]                               SLAVE_AWBURST;
  wire [NUM_SLAVES*2-1:0]                               SLAVE_AWLOCK;
  wire [NUM_SLAVES*4-1:0]                               SLAVE_AWCACHE;
  wire [NUM_SLAVES*3-1:0]                               SLAVE_AWPROT;
  wire [NUM_SLAVES*4-1:0]                               SLAVE_AWREGION;
  wire [NUM_SLAVES*4-1:0]                               SLAVE_AWQOS;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                      SLAVE_AWUSER;
  wire [NUM_SLAVES-1:0]                                 SLAVE_AWVALID;
  wire [NUM_SLAVES-1:0]                                 SLAVE_AWREADY;
  
  //====================== Slave Write Data Ports  ====================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE_WID;
  wire [SLAVE_DATA_WIDTH_PORT-1:0]                      SLAVE_WDATA;
  wire [SLAVE_DATA_WIDTH_PORT/8-1:0]                    SLAVE_WSTRB;
  wire [NUM_SLAVES-1:0]                                 SLAVE_WLAST;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                      SLAVE_WUSER;
  wire [NUM_SLAVES-1:0]                                 SLAVE_WVALID;
  wire [NUM_SLAVES-1:0]                                 SLAVE_WREADY;

  //====================== Slave Write Response Ports  ====================================================//
  wire [NUM_SLAVES*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0]    SLAVE_BID;
  wire [NUM_SLAVES*2-1:0]                               SLAVE_BRESP;
  wire [NUM_SLAVES*USER_WIDTH-1:0]                      SLAVE_BUSER;
  wire [NUM_SLAVES-1:0]                                 SLAVE_BVALID;
  wire [NUM_SLAVES-1:0]                                 SLAVE_BREADY;
       
  //====================== Master Read Address Ports  ================================================//
  wire [NUM_MASTERS*ID_WIDTH-1:0]                       masterARID;
  wire [NUM_MASTERS*ADDR_WIDTH-1:0]                     masterARADDR;
  wire [NUM_MASTERS*8-1:0]                              masterARLEN;
  wire [NUM_MASTERS*3-1:0]                              masterARSIZE;
  wire [NUM_MASTERS*2-1:0]                              masterARBURST;
  wire [NUM_MASTERS*2-1:0]                              masterARLOCK;
  wire [NUM_MASTERS*4-1:0]                              masterARCACHE;
  wire [NUM_MASTERS*3-1:0]                              masterARPROT;
  wire [NUM_MASTERS*4-1:0]                              masterARREGION;
  wire [NUM_MASTERS*4-1:0]                              masterARQOS;    // not used
  wire [NUM_MASTERS*USER_WIDTH-1:0]                     masterARUSER;
  wire [NUM_MASTERS-1:0]                                masterARVALID;
  wire [NUM_MASTERS-1:0]                                masterARREADY;
    
  //====================== Master Read Data Ports  ===================================================//
  wire [NUM_MASTERS*ID_WIDTH-1:0]                       masterRID;
  wire [NUM_MASTERS*DATA_WIDTH-1:0]                     masterRDATA;
  wire [NUM_MASTERS*2-1:0]                              masterRRESP;
  wire [NUM_MASTERS-1:0]                                masterRLAST;
  wire [NUM_MASTERS*USER_WIDTH-1:0]                     masterRUSER;
  wire [NUM_MASTERS-1:0]                                masterRVALID;

  wire [NUM_MASTERS-1:0]                                masterRREADY;
   
  //====================== Master Write Address Ports  ===================================================//
  wire [NUM_MASTERS*ID_WIDTH-1:0]                       masterAWID;
  wire [NUM_MASTERS*ADDR_WIDTH-1:0]                     masterAWADDR;
  wire [NUM_MASTERS*8-1:0]                              masterAWLEN;
  wire [NUM_MASTERS*3-1:0]                              masterAWSIZE;
  wire [NUM_MASTERS*2-1:0]                              masterAWBURST;
  wire [NUM_MASTERS*2-1:0]                              masterAWLOCK;
  wire [NUM_MASTERS*4-1:0]                              masterAWCACHE;
  wire [NUM_MASTERS*3-1:0]                              masterAWPROT;
  wire [NUM_MASTERS*4-1:0]                              masterAWREGION;
  wire [NUM_MASTERS*4-1:0]                              masterAWQOS;        // not used
  wire [NUM_MASTERS*USER_WIDTH-1:0]                     masterAWUSER;        // not used
  wire [NUM_MASTERS-1:0]                                masterAWVALID;
  wire [NUM_MASTERS-1:0]                                masterAWREADY;
    
  //====================== Master Write Data Ports  ===================================================//
  wire [NUM_MASTERS*DATA_WIDTH-1:0]                     masterWDATA;
  wire [NUM_MASTERS*DATA_WIDTH/8-1:0]                   masterWSTRB;
  wire [NUM_MASTERS-1:0]                                masterWLAST;
  wire [NUM_MASTERS*USER_WIDTH-1:0]                     masterWUSER;
  wire [NUM_MASTERS-1:0]                                masterWVALID;
  wire [NUM_MASTERS-1:0]                                masterWREADY;
 
  //====================== Master Write Response Ports  ===================================================//
  wire [NUM_MASTERS*ID_WIDTH-1:0]                       masterBID;
  wire [NUM_MASTERS*2-1:0]                              masterBRESP;
  wire [NUM_MASTERS*USER_WIDTH-1:0]                     masterBUSER;
  wire [NUM_MASTERS-1:0]                                masterBVALID;
  wire [NUM_MASTERS-1:0]                                masterBREADY;



  //==============================Wires between Master inputs/outputs And caxi4interconnect_MasterConvertor=============================
  // CB Master Write Address Ports
  wire [NUM_MASTERS*ID_WIDTH-1:0]                     MASTER_AWID;
  wire [NUM_MASTERS*ADDR_WIDTH-1:0]                   MASTER_AWADDR;
  wire [NUM_MASTERS*8-1:0]                            MASTER_AWLEN;
  wire [NUM_MASTERS*3-1:0]                            MASTER_AWSIZE;
  wire [NUM_MASTERS*2-1:0]                            MASTER_AWBURST;
  wire [NUM_MASTERS*2-1:0]                            MASTER_AWLOCK;
  wire [NUM_MASTERS*4-1:0]                            MASTER_AWCACHE;
  wire [NUM_MASTERS*3-1:0]                            MASTER_AWPROT;
  wire [NUM_MASTERS*4-1:0]                            MASTER_AWQOS;      // not used
  wire [NUM_MASTERS*USER_WIDTH-1:0]                   MASTER_AWUSER;      // not used
  wire [NUM_MASTERS-1:0]                              MASTER_AWVALID;
  wire [NUM_MASTERS-1:0]                              MASTER_AWREADY;
  wire [NUM_MASTERS*4-1:0]                            MASTER_AWREGION;
  
  // CB Master Write Data Ports
  wire [MASTER_DATA_WIDTH_PORT-1:0]                   MASTER_WDATA;
  wire [MASTER_DATA_WIDTH_PORT/8-1:0]                 MASTER_WSTRB;
  wire [NUM_MASTERS-1:0]                              MASTER_WLAST;
  wire [NUM_MASTERS*USER_WIDTH-1:0]                   MASTER_WUSER;
  wire [NUM_MASTERS-1:0]                              MASTER_WVALID;
  wire [NUM_MASTERS-1:0]                              MASTER_WREADY;
                                              
  // CB Master Write Response Ports
  wire [NUM_MASTERS*ID_WIDTH-1:0]                     MASTER_BID;
  wire [NUM_MASTERS*2-1:0]                            MASTER_BRESP;
  wire [NUM_MASTERS*USER_WIDTH-1:0]                   MASTER_BUSER;
  wire [NUM_MASTERS-1:0]                              MASTER_BVALID;
  wire [NUM_MASTERS-1:0]                              MASTER_BREADY;

  // CB Master Read Address Ports
  wire [NUM_MASTERS*ID_WIDTH-1:0]                     MASTER_ARID;
  wire [NUM_MASTERS*ADDR_WIDTH-1:0]                   MASTER_ARADDR;
  wire [NUM_MASTERS*8-1:0]                            MASTER_ARLEN;
  wire [NUM_MASTERS*3-1:0]                            MASTER_ARSIZE;
  wire [NUM_MASTERS*2-1:0]                            MASTER_ARBURST;
  wire [NUM_MASTERS*2-1:0]                            MASTER_ARLOCK;
  wire [NUM_MASTERS*4-1:0]                            MASTER_ARCACHE;
  wire [NUM_MASTERS*3-1:0]                            MASTER_ARPROT;
  wire [NUM_MASTERS*4-1:0]                            MASTER_ARREGION;
  wire [NUM_MASTERS*4-1:0]                            MASTER_ARQOS;    // not used
  wire [NUM_MASTERS*USER_WIDTH-1:0]                   MASTER_ARUSER;
  wire [NUM_MASTERS-1:0]                              MASTER_ARVALID;
  wire [NUM_MASTERS-1:0]                              MASTER_ARREADY;

  // CB Master Read Data Ports
  wire [NUM_MASTERS*ID_WIDTH-1:0]                     MASTER_RID;
  wire [MASTER_DATA_WIDTH_PORT-1:0]                   MASTER_RDATA;
  wire [NUM_MASTERS*2-1:0]                            MASTER_RRESP;
  wire [NUM_MASTERS-1:0]                              MASTER_RLAST;
  wire [NUM_MASTERS*USER_WIDTH-1:0]                   MASTER_RUSER;
  wire [NUM_MASTERS-1:0]                              MASTER_RVALID;
  wire [NUM_MASTERS-1:0]                              MASTER_RREADY;

        // AHB interface
  wire[8*32-1:0]                                      MASTER_HADDR;
  wire[8*3-1:0]                                       MASTER_HBURST;
  wire[7:0]                                           MASTER_HMASTLOCK;
  wire[8*7-1:0]                                       MASTER_HPROT;          
  wire[8*3-1:0]                                       MASTER_HSIZE;
  wire[7:0]                                           MASTER_HNONSEC;
  wire[8*2:0]                                         MASTER_HTRANS;
  wire[MASTER_DATA_WIDTH_PORT-1:0]                    MASTER_HWDATA;
  wire[MASTER_DATA_WIDTH_PORT-1:0]                    MASTER_HRDATA;
  wire[7:0]                                           MASTER_HWRITE;
  wire[7:0]                                           MASTER_HREADY;
  wire[7:0]                                           MASTER_HRESP;
  // wire[7:0]                                           MASTER_HEXOKAY;
  // wire[7:0]                                           MASTER_HEXCL;
  wire[7:0]                                           MASTER_HSEL;

  wire[8-1:0] M_CLK;
  wire[32-1:0] S_CLK;

   //SAR77215 fix
  //========================== Wire declarations for modified master QoS and Region signals ================ 
   

  wire [3:0]      MOD_MASTER0_AWREGION,  MOD_MASTER1_AWREGION,  MOD_MASTER2_AWREGION,  MOD_MASTER3_AWREGION,  MOD_MASTER4_AWREGION,  MOD_MASTER5_AWREGION,  MOD_MASTER6_AWREGION,  MOD_MASTER7_AWREGION;
  wire [3:0]      MOD_MASTER0_AWQOS,     MOD_MASTER1_AWQOS,     MOD_MASTER2_AWQOS,     MOD_MASTER3_AWQOS,     MOD_MASTER4_AWQOS,     MOD_MASTER5_AWQOS,     MOD_MASTER6_AWQOS,     MOD_MASTER7_AWQOS;
  wire [3:0]      MOD_MASTER0_ARREGION,  MOD_MASTER1_ARREGION,  MOD_MASTER2_ARREGION,  MOD_MASTER3_ARREGION,  MOD_MASTER4_ARREGION,  MOD_MASTER5_ARREGION,  MOD_MASTER6_ARREGION,  MOD_MASTER7_ARREGION;
  wire [3:0]      MOD_MASTER0_ARQOS,     MOD_MASTER1_ARQOS,     MOD_MASTER2_ARQOS,     MOD_MASTER3_ARQOS,     MOD_MASTER4_ARQOS,     MOD_MASTER5_ARQOS,     MOD_MASTER6_ARQOS,     MOD_MASTER7_ARQOS;   
  
  //=========================== Wire declarations for ARESETN synchronizer in ACLK domain ==================
  
  wire            ACLK_syncReset;
   
   //========================== Zero Master Region and QoS values fir master type 3  (AXI3) (tc:) ===========
   
  assign  MOD_MASTER0_AWQOS    = (MASTER0_TYPE == 2'b11) ? 4'b0 : MASTER0_AWQOS;
  assign  MOD_MASTER0_AWREGION = (MASTER0_TYPE == 2'b11) ? 4'b0 : MASTER0_AWREGION;
  assign  MOD_MASTER0_ARQOS    = (MASTER0_TYPE == 2'b11) ? 4'b0 : MASTER0_ARQOS;
  assign  MOD_MASTER0_ARREGION = (MASTER0_TYPE == 2'b11) ? 4'b0 : MASTER0_ARREGION;
   
  assign  MOD_MASTER1_AWQOS    = (MASTER1_TYPE == 2'b11) ? 4'b0 : MASTER1_AWQOS;
  assign  MOD_MASTER1_AWREGION = (MASTER1_TYPE == 2'b11) ? 4'b0 : MASTER1_AWREGION;
  assign  MOD_MASTER1_ARQOS    = (MASTER1_TYPE == 2'b11) ? 4'b0 : MASTER1_ARQOS;
  assign  MOD_MASTER1_ARREGION = (MASTER1_TYPE == 2'b11) ? 4'b0 : MASTER1_ARREGION;
   
  assign  MOD_MASTER2_AWQOS    = (MASTER2_TYPE == 2'b11) ? 4'b0 : MASTER2_AWQOS;
  assign  MOD_MASTER2_AWREGION = (MASTER2_TYPE == 2'b11) ? 4'b0 : MASTER2_AWREGION;
  assign  MOD_MASTER2_ARQOS    = (MASTER2_TYPE == 2'b11) ? 4'b0 : MASTER2_ARQOS;
  assign  MOD_MASTER2_ARREGION = (MASTER2_TYPE == 2'b11) ? 4'b0 : MASTER2_ARREGION;

  assign  MOD_MASTER3_AWQOS    = (MASTER3_TYPE == 2'b11) ? 4'b0 : MASTER3_AWQOS;
  assign  MOD_MASTER3_AWREGION = (MASTER3_TYPE == 2'b11) ? 4'b0 : MASTER3_AWREGION;
  assign  MOD_MASTER3_ARQOS    = (MASTER3_TYPE == 2'b11) ? 4'b0 : MASTER3_ARQOS;
  assign  MOD_MASTER3_ARREGION = (MASTER3_TYPE == 2'b11) ? 4'b0 : MASTER3_ARREGION;
  
  assign  MOD_MASTER4_AWQOS    = (MASTER4_TYPE == 2'b11) ? 4'b0 : MASTER4_AWQOS;
  assign  MOD_MASTER4_AWREGION = (MASTER4_TYPE == 2'b11) ? 4'b0 : MASTER4_AWREGION;
  assign  MOD_MASTER4_ARQOS    = (MASTER4_TYPE == 2'b11) ? 4'b0 : MASTER4_ARQOS;
  assign  MOD_MASTER4_ARREGION = (MASTER4_TYPE == 2'b11) ? 4'b0 : MASTER4_ARREGION;
   
  assign  MOD_MASTER5_AWQOS    = (MASTER5_TYPE == 2'b11) ? 4'b0 : MASTER5_AWQOS;
  assign  MOD_MASTER5_AWREGION = (MASTER5_TYPE == 2'b11) ? 4'b0 : MASTER5_AWREGION;
  assign  MOD_MASTER5_ARQOS    = (MASTER5_TYPE == 2'b11) ? 4'b0 : MASTER5_ARQOS;
  assign  MOD_MASTER5_ARREGION = (MASTER5_TYPE == 2'b11) ? 4'b0 : MASTER5_ARREGION;
   
  assign  MOD_MASTER6_AWQOS    = (MASTER6_TYPE == 2'b11) ? 4'b0 : MASTER6_AWQOS;
  assign  MOD_MASTER6_AWREGION = (MASTER6_TYPE == 2'b11) ? 4'b0 : MASTER6_AWREGION;
  assign  MOD_MASTER6_ARQOS    = (MASTER6_TYPE == 2'b11) ? 4'b0 : MASTER6_ARQOS;
  assign  MOD_MASTER6_ARREGION = (MASTER6_TYPE == 2'b11) ? 4'b0 : MASTER6_ARREGION;
   
  assign  MOD_MASTER7_AWQOS    = (MASTER7_TYPE == 2'b11) ? 4'b0 : MASTER7_AWQOS;
  assign  MOD_MASTER7_AWREGION = (MASTER7_TYPE == 2'b11) ? 4'b0 : MASTER7_AWREGION;
  assign  MOD_MASTER7_ARQOS    = (MASTER7_TYPE == 2'b11) ? 4'b0 : MASTER7_ARQOS;
  assign  MOD_MASTER7_ARREGION = (MASTER7_TYPE == 2'b11) ? 4'b0 : MASTER7_ARREGION;
    
  //==============================Master Combine Signals===============================================

  //===================================================================================================
  // MASTER 0
  //===================================================================================================

  //output to master converter   

  assign  MASTER_ARID[(0+1)*ID_WIDTH-1:0*ID_WIDTH]                                        = MASTER0_ARID;
  assign  MASTER_ARADDR[(0+1)*ADDR_WIDTH-1:0*ADDR_WIDTH]                                  = MASTER0_ARADDR;
  assign  MASTER_ARLEN[(0+1)*8-1:0*8]                                                     = MASTER0_ARLEN;
  assign  MASTER_ARSIZE[(0+1)*3-1:0*3]                                                    = MASTER0_ARSIZE;
  assign  MASTER_ARBURST[(0+1)*2-1:0*2]                                                   = MASTER0_ARBURST;
  assign  MASTER_ARLOCK[(0+1)*2-1:0*2]                                                    = MASTER0_ARLOCK;
  assign  MASTER_ARCACHE[(0+1)*4-1:0*4]                                                   = MASTER0_ARCACHE;
  assign  MASTER_ARPROT[(0+1)*3-1:0*3]                                                    = MASTER0_ARPROT;
  assign  MASTER_ARREGION[(0+1)*4-1:0*4]                                                  = MOD_MASTER0_ARREGION;
  assign  MASTER_ARQOS[(0+1)*4-1:0*4]                                                     = MOD_MASTER0_ARQOS;
  assign  MASTER_ARUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH]                                  = MASTER0_ARUSER;
  assign  MASTER_ARVALID[0]                                                               = MASTER0_ARVALID;
  assign  MASTER_AWQOS[(0+1)*4-1:0*4]                                                     = MOD_MASTER0_AWQOS;
  assign  MASTER_AWREGION[(0+1)*4-1:0*4]                                                  = MOD_MASTER0_AWREGION;
  assign  MASTER_AWID[(0+1)*ID_WIDTH-1:0*ID_WIDTH]                                        = MASTER0_AWID;  
  assign  MASTER_AWADDR[(0+1)*ADDR_WIDTH-1:0*ADDR_WIDTH]                                  = MASTER0_AWADDR;  
  assign  MASTER_AWLEN[(0+1)*8-1:0*8]                                                     = MASTER0_AWLEN;  
  assign  MASTER_AWSIZE[(0+1)*3-1:0*3]                                                    = MASTER0_AWSIZE;  
  assign  MASTER_AWBURST[(0+1)*2-1:0*2]                                                   = MASTER0_AWBURST;  
  assign  MASTER_AWLOCK[(0+1)*2-1:0*2]                                                    = MASTER0_AWLOCK;  
  assign  MASTER_AWCACHE[(0+1)*4-1:0*4]                                                   = MASTER0_AWCACHE;  
  assign  MASTER_AWPROT[(0+1)*3-1:0*3]                                                    = MASTER0_AWPROT;  
  assign  MASTER_AWUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH]                                  = MASTER0_AWUSER;  
  assign  MASTER_AWVALID[0]                                                               = MASTER0_AWVALID;  
  assign  MASTER_WDATA[MDW_UPPER_VEC[(0+1)*13-1:13*0]-1:MDW_LOWER_VEC[(0+1)*13-1:13*0]]   = MASTER0_WDATA;  
  assign  MASTER_WSTRB[MDW_UPPER_VEC[(0+1)*13-1:13*0]/8-1:MDW_LOWER_VEC[(0+1)*13-1:13*0]] = MASTER0_WSTRB;  
  assign  MASTER_WLAST[0]                                                                 = MASTER0_WLAST;  
  assign  MASTER_WUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH]                                   = MASTER0_WUSER;  
  assign  MASTER_WVALID[0]                                                                = MASTER0_WVALID;  
  assign  MASTER_BREADY[0]                                                                = MASTER0_BREADY;  
  assign  MASTER_RREADY[0]                                                                = MASTER0_RREADY;

  assign  MASTER0_RID           = MASTER_RID[(0+1)*ID_WIDTH-1:0*ID_WIDTH];
  assign  MASTER0_RDATA         = MASTER_RDATA[MDW_UPPER_VEC[(0+1)*13-1:13*0]-1:MDW_LOWER_VEC[(0+1)*13-1:13*0]];
  assign  MASTER0_RRESP         = MASTER_RRESP[(0+1)*2-1:0*2];
  assign  MASTER0_RUSER         = MASTER_RUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH];
  assign  MASTER0_BID           = MASTER_BID[(0+1)*ID_WIDTH-1:0*ID_WIDTH];
  assign  MASTER0_BRESP         = MASTER_BRESP[(0+1)*2-1:0*2];
  assign  MASTER0_BUSER         = MASTER_BUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH];
  assign  MASTER0_ARREADY       = MASTER_ARREADY[0];
  assign  MASTER0_RLAST         = MASTER_RLAST[0];
  assign  MASTER0_RVALID        = MASTER_RVALID[0];
  assign  MASTER0_AWREADY       = MASTER_AWREADY[0];
  assign  MASTER0_WREADY        = MASTER_WREADY[0];
  assign  MASTER0_BVALID        = MASTER_BVALID[0];

        // AHB interface
  assign MASTER_HADDR[32*(0+1)-1:32*0]                                                    = MASTER0_HADDR;
  assign MASTER_HBURST[3*(0+1)-1:3*0]                                                     = MASTER0_HBURST;
  assign MASTER_HMASTLOCK[0]                                                              = MASTER0_HMASTLOCK;
  assign MASTER_HPROT[7*(0+1)-1:7*0]                                                      = MASTER0_HPROT;          
  assign MASTER_HSIZE[3*(0+1)-1:3*0]                                                      = MASTER0_HSIZE;
  assign MASTER_HNONSEC[0]                                                                = MASTER0_HNONSEC;
  assign MASTER_HTRANS[2*(0+1)-1:2*0]                                                     = MASTER0_HTRANS;
  assign MASTER_HWDATA[MDW_UPPER_VEC[(0+1)*13-1:13*0]-1:MDW_LOWER_VEC[(0+1)*13-1:13*0]]   = MASTER0_HWDATA;
  assign MASTER0_HRDATA                                                                   = MASTER_HRDATA[MDW_UPPER_VEC[(0+1)*13-1:13*0]-1:MDW_LOWER_VEC[(0+1)*13-1:13*0]];
  assign MASTER_HWRITE[0]                                                                 = MASTER0_HWRITE;
  assign MASTER0_HRESP                                                                    = MASTER_HRESP[0];
  // assign MASTER0_HEXOKAY                                                                  = MASTER_HEXOKAY[0];
  // assign MASTER_HEXCL[0]                                                                  = MASTER0_HEXCL;
  assign MASTER_HSEL[0]                                                                   = MASTER0_HSEL;
  assign MASTER0_HREADY                                                                   = MASTER_HREADY[0];

  //===================================================================================================
  //MASTER 1
  //===================================================================================================  

  if ( NUM_MASTERS > 1)
    begin
      //output to master converter 
      
      assign   MASTER_ARID[(1+1)*ID_WIDTH-1:1*ID_WIDTH]                                         = MASTER1_ARID;
      assign   MASTER_ARADDR[(1+1)*ADDR_WIDTH-1:1*ADDR_WIDTH]                                   = MASTER1_ARADDR;
      assign   MASTER_ARLEN[(1+1)*8-1:1*8]                                                      = MASTER1_ARLEN;
      assign   MASTER_ARSIZE[(1+1)*3-1:1*3]                                                     = MASTER1_ARSIZE;
      assign   MASTER_ARBURST[(1+1)*2-1:1*2]                                                    = MASTER1_ARBURST;
      assign   MASTER_ARLOCK[(1+1)*2-1:1*2]                                                     = MASTER1_ARLOCK;
      assign   MASTER_ARCACHE[(1+1)*4-1:1*4]                                                    = MASTER1_ARCACHE;
      assign   MASTER_ARPROT[(1+1)*3-1:1*3]                                                     = MASTER1_ARPROT;
      assign   MASTER_ARREGION[(1+1)*4-1:1*4]                                                   = MOD_MASTER1_ARREGION;
      assign   MASTER_ARQOS[(1+1)*4-1:1*4]                                                      = MOD_MASTER1_ARQOS;
      assign   MASTER_ARUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH]                                   = MASTER1_ARUSER;
      assign   MASTER_ARVALID[1]                                                                = MASTER1_ARVALID;
      assign   MASTER_AWQOS[(1+1)*4-1:1*4]                                                      = MOD_MASTER1_AWQOS;
      assign   MASTER_AWREGION[(1+1)*4-1:1*4]                                                   = MOD_MASTER1_AWREGION;
      assign  MASTER_AWID[(1+1)*ID_WIDTH-1:1*ID_WIDTH]                                          = MASTER1_AWID;  
      assign  MASTER_AWADDR[(1+1)*ADDR_WIDTH-1:1*ADDR_WIDTH]                                    = MASTER1_AWADDR;  
      assign  MASTER_AWLEN[(1+1)*8-1:1*8]                                                       = MASTER1_AWLEN;  
      assign  MASTER_AWSIZE[(1+1)*3-1:1*3]                                                      = MASTER1_AWSIZE;  
      assign  MASTER_AWBURST[(1+1)*2-1:1*2]                                                     = MASTER1_AWBURST;  
      assign  MASTER_AWLOCK[(1+1)*2-1:1*2]                                                      = MASTER1_AWLOCK;  
      assign  MASTER_AWCACHE[(1+1)*4-1:1*4]                                                     = MASTER1_AWCACHE;  
      assign  MASTER_AWPROT[(1+1)*3-1:1*3]                                                      = MASTER1_AWPROT;  
      assign  MASTER_AWUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH]                                    = MASTER1_AWUSER;  
      assign  MASTER_AWVALID[1]                                                                 = MASTER1_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(1+1)*13-1:13*1]-1:MDW_LOWER_VEC[(1+1)*13-1:13*1]]     = MASTER1_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(1+1)*13-1:13*1]/8-1:MDW_LOWER_VEC[(1+1)*13-1:13*1]/8] = MASTER1_WSTRB;  
      assign  MASTER_WLAST[1]                                                                   = MASTER1_WLAST;  
      assign  MASTER_WUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH]                                     = MASTER1_WUSER;  
      assign  MASTER_WVALID[1]                                                                  = MASTER1_WVALID;  
      assign  MASTER_BREADY[1]                                                                  = MASTER1_BREADY;  
      assign  MASTER_RREADY[1]                                                                  = MASTER1_RREADY;  

      assign MASTER1_RID        = MASTER_RID[(1+1)*ID_WIDTH-1:1*ID_WIDTH];
      assign MASTER1_RDATA      = MASTER_RDATA[MDW_UPPER_VEC[(1+1)*13-1:13*1]-1:MDW_LOWER_VEC[(1+1)*13-1:13*1]];
      assign MASTER1_RRESP      = MASTER_RRESP[(1+1)*2-1:1*2];
      assign MASTER1_RUSER      = MASTER_RUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH];
      assign MASTER1_BID        = MASTER_BID[(1+1)*ID_WIDTH-1:1*ID_WIDTH];
      assign MASTER1_BRESP      = MASTER_BRESP[(1+1)*2-1:1*2];
      assign MASTER1_BUSER      = MASTER_BUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH];
      assign MASTER1_ARREADY    = MASTER_ARREADY[1];
      assign MASTER1_RLAST      = MASTER_RLAST[1];
      assign MASTER1_RVALID     = MASTER_RVALID[1];
      assign MASTER1_AWREADY    = MASTER_AWREADY[1];
      assign MASTER1_WREADY     = MASTER_WREADY[1];
      assign MASTER1_BVALID     = MASTER_BVALID[1];

      // AHB interface
      assign MASTER_HADDR[32*(1+1)-1:32*1]                                                  = MASTER1_HADDR;
      assign MASTER_HBURST[3*(1+1)-1:3*1]                                                   = MASTER1_HBURST;
      assign MASTER_HMASTLOCK[1]                                                            = MASTER1_HMASTLOCK;
      assign MASTER_HPROT[7*(1+1)-1:7*1]                                                    = MASTER1_HPROT;          
      assign MASTER_HSIZE[3*(1+1)-1:3*1]                                                    = MASTER1_HSIZE;
      assign MASTER_HNONSEC[1]                                                              = MASTER1_HNONSEC;
      assign MASTER_HTRANS[2*(1+1)-1:2*1]                                                   = MASTER1_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(1+1)*13-1:13*1]-1:MDW_LOWER_VEC[(1+1)*13-1:13*1]] = MASTER1_HWDATA;
      assign MASTER1_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(1+1)*13-1:13*1]-1:MDW_LOWER_VEC[(1+1)*13-1:13*1]];
      assign MASTER_HWRITE[1]                                                               = MASTER1_HWRITE;
      assign MASTER1_HRESP                                                                  = MASTER_HRESP[1];
//      assign MASTER1_HEXOKAY                                                              = MASTER_HEXOKAY[1];
//    assign MASTER_HEXCL[1]                                                                = MASTER1_HEXCL;
      assign MASTER_HSEL[1]                                                                 = MASTER1_HSEL;
      assign MASTER1_HREADY                                                                 = MASTER_HREADY[1];

    end

  //===================================================================================================
  //MASTER 2
  //===================================================================================================
  if ( NUM_MASTERS > 2 )
    begin
      //output to master converter 
      assign  MASTER_ARID[(2+1)*ID_WIDTH-1:2*ID_WIDTH]                                          = MASTER2_ARID;
      assign  MASTER_ARADDR[(2+1)*ADDR_WIDTH-1:2*ADDR_WIDTH]                                    = MASTER2_ARADDR;
      assign  MASTER_ARLEN[(2+1)*8-1:2*8]                                                       = MASTER2_ARLEN;
      assign  MASTER_ARSIZE[(2+1)*3-1:2*3]                                                      = MASTER2_ARSIZE;
      assign  MASTER_ARBURST[(2+1)*2-1:2*2]                                                     = MASTER2_ARBURST;
      assign  MASTER_ARLOCK[(2+1)*2-1:2*2]                                                      = MASTER2_ARLOCK;
      assign  MASTER_ARCACHE[(2+1)*4-1:2*4]                                                     = MASTER2_ARCACHE;
      assign  MASTER_ARPROT[(2+1)*3-1:2*3]                                                      = MASTER2_ARPROT;
      assign  MASTER_ARREGION[(2+1)*4-1:2*4]                                                    = MOD_MASTER2_ARREGION;
      assign  MASTER_ARQOS[(2+1)*4-1:2*4]                                                       = MOD_MASTER2_ARQOS;
      assign  MASTER_ARUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH]                                    = MASTER2_ARUSER;
      assign  MASTER_ARVALID[2]                                                                 = MASTER2_ARVALID;
      assign  MASTER_AWQOS[(2+1)*4-1:2*4]                                                       = MOD_MASTER2_AWQOS;
      assign  MASTER_AWREGION[(2+1)*4-1:2*4]                                                    = MOD_MASTER2_AWREGION;
      assign  MASTER_AWID[(2+1)*ID_WIDTH-1:2*ID_WIDTH]                                          = MASTER2_AWID;  
      assign  MASTER_AWADDR[(2+1)*ADDR_WIDTH-1:2*ADDR_WIDTH]                                    = MASTER2_AWADDR;  
      assign  MASTER_AWLEN[(2+1)*8-1:2*8]                                                       = MASTER2_AWLEN;  
      assign  MASTER_AWSIZE[(2+1)*3-1:2*3]                                                      = MASTER2_AWSIZE;  
      assign  MASTER_AWBURST[(2+1)*2-1:2*2]                                                     = MASTER2_AWBURST;  
      assign  MASTER_AWLOCK[(2+1)*2-1:2*2]                                                      = MASTER2_AWLOCK;  
      assign  MASTER_AWCACHE[(2+1)*4-1:2*4]                                                     = MASTER2_AWCACHE;  
      assign  MASTER_AWPROT[(2+1)*3-1:2*3]                                                      = MASTER2_AWPROT;  
      assign  MASTER_AWUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH]                                    = MASTER2_AWUSER;  
      assign  MASTER_AWVALID[2]                                                                 = MASTER2_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(2+1)*13-1:13*2]-1:MDW_LOWER_VEC[(2+1)*13-1:13*2]]     = MASTER2_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(2+1)*13-1:13*2]/8-1:MDW_LOWER_VEC[(2+1)*13-1:13*2]/8] = MASTER2_WSTRB;  
      assign  MASTER_WLAST[2]                                                                   = MASTER2_WLAST;  
      assign  MASTER_WUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH]                                     = MASTER2_WUSER;  
      assign  MASTER_WVALID[2]                                                                  = MASTER2_WVALID;  
      assign  MASTER_BREADY[2]                                                                  = MASTER2_BREADY;  
      assign  MASTER_RREADY[2]                                                                  = MASTER2_RREADY;  

      assign MASTER2_RID        = MASTER_RID[(2+1)*ID_WIDTH-1:2*ID_WIDTH];
      assign MASTER2_RDATA      = MASTER_RDATA[MDW_UPPER_VEC[(2+1)*13-1:13*2]-1:MDW_LOWER_VEC[(2+1)*13-1:13*2]];
      assign MASTER2_RRESP      = MASTER_RRESP[(2+1)*2-1:2*2];
      assign MASTER2_RUSER      = MASTER_RUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH];
      assign MASTER2_BID        = MASTER_BID[(2+1)*ID_WIDTH-1:2*ID_WIDTH];
      assign MASTER2_BRESP      = MASTER_BRESP[(2+1)*2-1:2*2];
      assign MASTER2_BUSER      = MASTER_BUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH];
      assign MASTER2_ARREADY    = MASTER_ARREADY[2];
      assign MASTER2_RLAST      = MASTER_RLAST[2];
      assign MASTER2_RVALID     = MASTER_RVALID[2];
      assign MASTER2_AWREADY    = MASTER_AWREADY[2];
      assign MASTER2_WREADY     = MASTER_WREADY[2];
      assign MASTER2_BVALID     = MASTER_BVALID[2];

      // AHB interface
      assign MASTER_HADDR[32*(2+1)-1:32*2]                                                  = MASTER2_HADDR;
      assign MASTER_HBURST[3*(2+1)-1:3*2]                                                   = MASTER2_HBURST;
      assign MASTER_HMASTLOCK[2]                                                            = MASTER2_HMASTLOCK;
      assign MASTER_HPROT[7*(2+1)-1:7*2]                                                    = MASTER2_HPROT;          
      assign MASTER_HSIZE[3*(2+1)-1:3*2]                                                    = MASTER2_HSIZE;
      assign MASTER_HNONSEC[2]                                                              = MASTER2_HNONSEC;
      assign MASTER_HTRANS[2*(2+1)-1:2*2]                                                   = MASTER2_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(2+1)*13-1:13*2]-1:MDW_LOWER_VEC[(2+1)*13-1:13*2]] = MASTER2_HWDATA;
      assign MASTER2_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(2+1)*13-1:13*2]-1:MDW_LOWER_VEC[(2+1)*13-1:13*2]];
      assign MASTER_HWRITE[2]                                                               = MASTER2_HWRITE;
      assign MASTER2_HRESP                                                                  = MASTER_HRESP[2];
//      assign MASTER2_HEXOKAY                                                              = MASTER_HEXOKAY[2];
//                  assign MASTER_HEXCL[2]                                                  = MASTER2_HEXCL;
      assign MASTER_HSEL[2]                                                                 = MASTER2_HSEL;
      assign MASTER2_HREADY                                                                 = MASTER_HREADY[2];

    end
    
  //===================================================================================================
  // MASTER 3
  //===================================================================================================
  if ( NUM_MASTERS > 3)
    begin    
      //output to master converter 
      
      assign  MASTER_ARID[(3+1)*ID_WIDTH-1:3*ID_WIDTH]                                          = MASTER3_ARID;
      assign  MASTER_ARADDR[(3+1)*ADDR_WIDTH-1:3*ADDR_WIDTH]                                    = MASTER3_ARADDR;
      assign  MASTER_ARLEN[(3+1)*8-1:3*8]                                                       = MASTER3_ARLEN;
      assign  MASTER_ARSIZE[(3+1)*3-1:3*3]                                                      = MASTER3_ARSIZE;
      assign  MASTER_ARBURST[(3+1)*2-1:3*2]                                                     = MASTER3_ARBURST;
      assign  MASTER_ARLOCK[(3+1)*2-1:3*2]                                                      = MASTER3_ARLOCK;
      assign  MASTER_ARCACHE[(3+1)*4-1:3*4]                                                     = MASTER3_ARCACHE;
      assign  MASTER_ARPROT[(3+1)*3-1:3*3]                                                      = MASTER3_ARPROT;
      assign  MASTER_ARREGION[(3+1)*4-1:3*4]                                                    = MOD_MASTER3_ARREGION;
      assign  MASTER_ARQOS[(3+1)*4-1:3*4]                                                       = MOD_MASTER3_ARQOS;
      assign  MASTER_ARUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH]                                    = MASTER3_ARUSER;
      assign  MASTER_ARVALID[3]                                                                 = MASTER3_ARVALID;
      assign  MASTER_AWQOS[(3+1)*4-1:3*4]                                                       = MOD_MASTER3_AWQOS;
      assign  MASTER_AWREGION[(3+1)*4-1:3*4]                                                    = MOD_MASTER3_AWREGION;
      assign  MASTER_AWID[(3+1)*ID_WIDTH-1:3*ID_WIDTH]                                          = MASTER3_AWID;  
      assign  MASTER_AWADDR[(3+1)*ADDR_WIDTH-1:3*ADDR_WIDTH]                                    = MASTER3_AWADDR;  
      assign  MASTER_AWLEN[(3+1)*8-1:3*8]                                                       = MASTER3_AWLEN;  
      assign  MASTER_AWSIZE[(3+1)*3-1:3*3]                                                      = MASTER3_AWSIZE;  
      assign  MASTER_AWBURST[(3+1)*2-1:3*2]                                                     = MASTER3_AWBURST;  
      assign  MASTER_AWLOCK[(3+1)*2-1:3*2]                                                      = MASTER3_AWLOCK;  
      assign  MASTER_AWCACHE[(3+1)*4-1:3*4]                                                     = MASTER3_AWCACHE;  
      assign  MASTER_AWPROT[(3+1)*3-1:3*3]                                                      = MASTER3_AWPROT;  
      assign  MASTER_AWUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH]                                    = MASTER3_AWUSER;  
      assign  MASTER_AWVALID[3]                                                                 = MASTER3_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(3+1)*13-1:13*3]-1:MDW_LOWER_VEC[(3+1)*13-1:13*3]]     = MASTER3_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(3+1)*13-1:13*3]/8-1:MDW_LOWER_VEC[(3+1)*13-1:13*3]/8] = MASTER3_WSTRB;  
      assign  MASTER_WLAST[3]                                                                   = MASTER3_WLAST;  
      assign  MASTER_WUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH]                                     = MASTER3_WUSER;  
      assign  MASTER_WVALID[3]                                                                  = MASTER3_WVALID;  
      assign  MASTER_BREADY[3]                                                                  = MASTER3_BREADY;  
      assign  MASTER_RREADY[3]                                                                  = MASTER3_RREADY;  

      assign MASTER3_RID        = MASTER_RID[(3+1)*ID_WIDTH-1:3*ID_WIDTH];
      assign MASTER3_RDATA      = MASTER_RDATA[MDW_UPPER_VEC[(3+1)*13-1:13*3]-1:MDW_LOWER_VEC[(3+1)*13-1:13*3]];
      assign MASTER3_RRESP      = MASTER_RRESP[(3+1)*2-1:3*2];
      assign MASTER3_RUSER      = MASTER_RUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH];
      assign MASTER3_BID        = MASTER_BID[(3+1)*ID_WIDTH-1:3*ID_WIDTH];
      assign MASTER3_BRESP      = MASTER_BRESP[(3+1)*2-1:3*2];
      assign MASTER3_BUSER      = MASTER_BUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH];
      assign MASTER3_ARREADY    = MASTER_ARREADY[3];
      assign MASTER3_RLAST      = MASTER_RLAST[3];
      assign MASTER3_RVALID     = MASTER_RVALID[3];
      assign MASTER3_AWREADY    = MASTER_AWREADY[3];
      assign MASTER3_WREADY     = MASTER_WREADY[3];
      assign MASTER3_BVALID     = MASTER_BVALID[3];

      // AHB interface
      assign MASTER_HADDR[32*(3+1)-1:32*3]                                                  = MASTER3_HADDR;
      assign MASTER_HBURST[3*(3+1)-1:3*3]                                                   = MASTER3_HBURST;
      assign MASTER_HMASTLOCK[3]                                                            = MASTER3_HMASTLOCK;
      assign MASTER_HPROT[7*(3+1)-1:7*3]                                                    = MASTER3_HPROT;          
      assign MASTER_HSIZE[3*(3+1)-1:3*3]                                                    = MASTER3_HSIZE;
      assign MASTER_HNONSEC[3]                                                              = MASTER3_HNONSEC;
      assign MASTER_HTRANS[2*(3+1)-1:2*3]                                                   = MASTER3_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(3+1)*13-1:13*3]-1:MDW_LOWER_VEC[(3+1)*13-1:13*3]] = MASTER3_HWDATA;
      assign MASTER3_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(3+1)*13-1:13*3]-1:MDW_LOWER_VEC[(3+1)*13-1:13*3]];
      assign MASTER_HWRITE[3]                                                               = MASTER3_HWRITE;
      assign MASTER3_HRESP                                                                  = MASTER_HRESP[3];
//      assign MASTER3_HEXOKAY                                                              = MASTER_HEXOKAY[3];
//      assign MASTER_HEXCL[3]                                                              = MASTER3_HEXCL;
      assign MASTER_HSEL[3]                                                                 = MASTER3_HSEL;
      assign MASTER3_HREADY = MASTER_HREADY[3];
    end
    
  //===================================================================================================
  // MASTER 4
  //===================================================================================================
  if ( NUM_MASTERS > 4)
    begin  
      //output to master converter
      
      assign   MASTER_ARID[(4+1)*ID_WIDTH-1:4*ID_WIDTH]                                         = MASTER4_ARID;
      assign   MASTER_ARADDR[(4+1)*ADDR_WIDTH-1:4*ADDR_WIDTH]                                   = MASTER4_ARADDR;
      assign   MASTER_ARLEN[(4+1)*8-1:4*8]                                                      = MASTER4_ARLEN;
      assign   MASTER_ARSIZE[(4+1)*3-1:4*3]                                                     = MASTER4_ARSIZE;
      assign   MASTER_ARBURST[(4+1)*2-1:4*2]                                                    = MASTER4_ARBURST;
      assign   MASTER_ARLOCK[(4+1)*2-1:4*2]                                                     = MASTER4_ARLOCK;
      assign   MASTER_ARCACHE[(4+1)*4-1:4*4]                                                    = MASTER4_ARCACHE;
      assign   MASTER_ARPROT[(4+1)*3-1:4*3]                                                     = MASTER4_ARPROT;
      assign   MASTER_ARREGION[(4+1)*4-1:4*4]                                                   = MOD_MASTER4_ARREGION;
      assign   MASTER_ARQOS[(4+1)*4-1:4*4]                                                      = MOD_MASTER4_ARQOS;
      assign   MASTER_ARUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH]                                   = MASTER4_ARUSER;
      assign   MASTER_ARVALID[4]                                                                = MASTER4_ARVALID;
      assign   MASTER_AWQOS[(4+1)*4-1:4*4]                                                      = MOD_MASTER4_AWQOS;
      assign   MASTER_AWREGION[(4+1)*4-1:4*4]                                                   = MOD_MASTER4_AWREGION;
      assign  MASTER_AWID[(4+1)*ID_WIDTH-1:4*ID_WIDTH]                                          = MASTER4_AWID;  
      assign  MASTER_AWADDR[(4+1)*ADDR_WIDTH-1:4*ADDR_WIDTH]                                    = MASTER4_AWADDR;  
      assign  MASTER_AWLEN[(4+1)*8-1:4*8]                                                       = MASTER4_AWLEN;  
      assign  MASTER_AWSIZE[(4+1)*3-1:4*3]                                                      = MASTER4_AWSIZE;  
      assign  MASTER_AWBURST[(4+1)*2-1:4*2]                                                     = MASTER4_AWBURST;  
      assign  MASTER_AWLOCK[(4+1)*2-1:4*2]                                                      = MASTER4_AWLOCK;  
      assign  MASTER_AWCACHE[(4+1)*4-1:4*4]                                                     = MASTER4_AWCACHE;  
      assign  MASTER_AWPROT[(4+1)*3-1:4*3]                                                      = MASTER4_AWPROT;  
      assign  MASTER_AWUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH]                                    = MASTER4_AWUSER;  
      assign  MASTER_AWVALID[4]                                                                 = MASTER4_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(4+1)*13-1:13*4]-1:MDW_LOWER_VEC[(4+1)*13-1:13*4]]     = MASTER4_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(4+1)*13-1:13*4]/8-1:MDW_LOWER_VEC[(4+1)*13-1:13*4]/8] = MASTER4_WSTRB;  
      assign  MASTER_WLAST[4]                                                                   = MASTER4_WLAST;  
      assign  MASTER_WUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH]                                     = MASTER4_WUSER;  
      assign  MASTER_WVALID[4]                                                                  = MASTER4_WVALID;  
      assign  MASTER_BREADY[4]                                                                  = MASTER4_BREADY;  
      assign  MASTER_RREADY[4]                                                                  = MASTER4_RREADY;

      assign MASTER4_RID        = MASTER_RID[(4+1)*ID_WIDTH-1:4*ID_WIDTH];
      assign MASTER4_RDATA      = MASTER_RDATA[MDW_UPPER_VEC[(4+1)*13-1:13*4]-1:MDW_LOWER_VEC[(4+1)*13-1:13*4]];
      assign MASTER4_RRESP      = MASTER_RRESP[(4+1)*2-1:4*2];
      assign MASTER4_RUSER      = MASTER_RUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH];
      assign MASTER4_BID        = MASTER_BID[(4+1)*ID_WIDTH-1:4*ID_WIDTH];
      assign MASTER4_BRESP      = MASTER_BRESP[(4+1)*2-1:4*2];
      assign MASTER4_BUSER      = MASTER_BUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH];
      assign MASTER4_ARREADY    = MASTER_ARREADY[4];
      assign MASTER4_RLAST      = MASTER_RLAST[4];
      assign MASTER4_RVALID     = MASTER_RVALID[4];
      assign MASTER4_AWREADY    = MASTER_AWREADY[4];
      assign MASTER4_WREADY     = MASTER_WREADY[4];
      assign MASTER4_BVALID     = MASTER_BVALID[4];

      // AHB interface
      assign MASTER_HADDR[32*(4+1)-1:32*4]                                                  = MASTER4_HADDR;
      assign MASTER_HBURST[3*(4+1)-1:3*4]                                                   = MASTER4_HBURST;
      assign MASTER_HMASTLOCK[4]                                                            = MASTER4_HMASTLOCK;
      assign MASTER_HPROT[7*(4+1)-1:7*4]                                                    = MASTER4_HPROT;          
      assign MASTER_HSIZE[3*(4+1)-1:3*4]                                                    = MASTER4_HSIZE;
      assign MASTER_HNONSEC[4]                                                              = MASTER4_HNONSEC;
      assign MASTER_HTRANS[2*(4+1)-1:2*4]                                                   = MASTER4_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(4+1)*13-1:13*4]-1:MDW_LOWER_VEC[(4+1)*13-1:13*4]] = MASTER4_HWDATA;
      assign MASTER4_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(4+1)*13-1:13*4]-1:MDW_LOWER_VEC[(4+1)*13-1:13*4]];
      assign MASTER_HWRITE[4]                                                               = MASTER4_HWRITE;
      assign MASTER4_HRESP                                                                  = MASTER_HRESP[4];
//      assign MASTER4_HEXOKAY                                                              = MASTER_HEXOKAY[4];
//      assign MASTER_HEXCL[4]                                                              = MASTER4_HEXCL;
      assign MASTER_HSEL[4]                                                                 = MASTER4_HSEL;
      assign MASTER4_HREADY                                                                 = MASTER_HREADY[4];
    end
    
  //===================================================================================================
  // MASTER 5
  //===================================================================================================
  if ( NUM_MASTERS > 5)
    begin  
      //output to master converter 

      assign  MASTER_ARID[(5+1)*ID_WIDTH-1:5*ID_WIDTH]                                          = MASTER5_ARID;
      assign  MASTER_ARADDR[(5+1)*ADDR_WIDTH-1:5*ADDR_WIDTH]                                    = MASTER5_ARADDR;
      assign  MASTER_ARLEN[(5+1)*8-1:5*8]                                                       = MASTER5_ARLEN;
      assign  MASTER_ARSIZE[(5+1)*3-1:5*3]                                                      = MASTER5_ARSIZE;
      assign  MASTER_ARBURST[(5+1)*2-1:5*2]                                                     = MASTER5_ARBURST;
      assign  MASTER_ARLOCK[(5+1)*2-1:5*2]                                                      = MASTER5_ARLOCK;
      assign  MASTER_ARCACHE[(5+1)*4-1:5*4]                                                     = MASTER5_ARCACHE;
      assign  MASTER_ARPROT[(5+1)*3-1:5*3]                                                      = MASTER5_ARPROT;
      assign  MASTER_ARREGION[(5+1)*4-1:5*4]                                                    = MOD_MASTER5_ARREGION;
      assign  MASTER_ARQOS[(5+1)*4-1:5*4]                                                       = MOD_MASTER5_ARQOS;
      assign  MASTER_ARUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH]                                    = MASTER5_ARUSER;
      assign  MASTER_ARVALID[5]                                                                 = MASTER5_ARVALID;
      assign  MASTER_AWQOS[(5+1)*4-1:5*4]                                                       = MOD_MASTER5_AWQOS;
      assign  MASTER_AWREGION[(5+1)*4-1:5*4]                                                    = MOD_MASTER5_AWREGION;
      assign  MASTER_AWID[(5+1)*ID_WIDTH-1:5*ID_WIDTH]                                          = MASTER5_AWID;  
      assign  MASTER_AWADDR[(5+1)*ADDR_WIDTH-1:5*ADDR_WIDTH]                                    = MASTER5_AWADDR;  
      assign  MASTER_AWLEN[(5+1)*8-1:5*8]                                                       = MASTER5_AWLEN;  
      assign  MASTER_AWSIZE[(5+1)*3-1:5*3]                                                      = MASTER5_AWSIZE;  
      assign  MASTER_AWBURST[(5+1)*2-1:5*2]                                                     = MASTER5_AWBURST;  
      assign  MASTER_AWLOCK[(5+1)*2-1:5*2]                                                      = MASTER5_AWLOCK;  
      assign  MASTER_AWCACHE[(5+1)*4-1:5*4]                                                     = MASTER5_AWCACHE;  
      assign  MASTER_AWPROT[(5+1)*3-1:5*3]                                                      = MASTER5_AWPROT;  
      assign  MASTER_AWUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH]                                    = MASTER5_AWUSER;  
      assign  MASTER_AWVALID[5]                                                                 = MASTER5_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(5+1)*13-1:13*5]-1:MDW_LOWER_VEC[(5+1)*13-1:13*5]]     = MASTER5_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(5+1)*13-1:13*5]/8-1:MDW_LOWER_VEC[(5+1)*13-1:13*5]/8] = MASTER5_WSTRB;  
      assign  MASTER_WLAST[5]                                                                   = MASTER5_WLAST;  
      assign  MASTER_WUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH]                                     = MASTER5_WUSER;  
      assign  MASTER_WVALID[5]                                                                  = MASTER5_WVALID;  
      assign  MASTER_BREADY[5]                                                                  = MASTER5_BREADY;  
      assign  MASTER_RREADY[5]                                                                  = MASTER5_RREADY;

      assign  MASTER5_RID       = MASTER_RID[(5+1)*ID_WIDTH-1:5*ID_WIDTH];
      assign  MASTER5_RDATA     = MASTER_RDATA[MDW_UPPER_VEC[(5+1)*13-1:13*5]-1:MDW_LOWER_VEC[(5+1)*13-1:13*5]];
      assign  MASTER5_RRESP     = MASTER_RRESP[(5+1)*2-1:5*2];
      assign  MASTER5_RUSER     = MASTER_RUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH];
      assign  MASTER5_BID       = MASTER_BID[(5+1)*ID_WIDTH-1:5*ID_WIDTH];
      assign  MASTER5_BRESP     = MASTER_BRESP[(5+1)*2-1:5*2];
      assign  MASTER5_BUSER     = MASTER_BUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH];
      assign  MASTER5_ARREADY   = MASTER_ARREADY[5];
      assign  MASTER5_RLAST     = MASTER_RLAST[5];
      assign  MASTER5_RVALID    = MASTER_RVALID[5];
      assign  MASTER5_AWREADY   = MASTER_AWREADY[5];
      assign  MASTER5_WREADY    = MASTER_WREADY[5];
      assign  MASTER5_BVALID    = MASTER_BVALID[5];

      // AHB interface
      assign MASTER_HADDR[32*(5+1)-1:32*5]                                                  = MASTER5_HADDR;
      assign MASTER_HBURST[3*(5+1)-1:3*5]                                                   = MASTER5_HBURST;
      assign MASTER_HMASTLOCK[5]                                                            = MASTER5_HMASTLOCK;
      assign MASTER_HPROT[7*(5+1)-1:7*5]                                                    = MASTER5_HPROT;          
      assign MASTER_HSIZE[3*(5+1)-1:3*5]                                                    = MASTER5_HSIZE;
      assign MASTER_HNONSEC[5]                                                              = MASTER5_HNONSEC;
      assign MASTER_HTRANS[2*(5+1)-1:2*5]                                                   = MASTER5_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(5+1)*13-1:13*5]-1:MDW_LOWER_VEC[(5+1)*13-1:13*5]] = MASTER5_HWDATA;
      assign MASTER5_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(5+1)*13-1:13*5]-1:MDW_LOWER_VEC[(5+1)*13-1:13*5]];
      assign MASTER_HWRITE[5]                                                               = MASTER5_HWRITE;
      assign MASTER5_HRESP                                                                  = MASTER_HRESP[5];
//      assign MASTER5_HEXOKAY                                                              = MASTER_HEXOKAY[5];
//      assign MASTER_HEXCL[5]                                                              = MASTER5_HEXCL;
      assign MASTER_HSEL[5]                                                                 = MASTER5_HSEL;
      assign MASTER5_HREADY                                                                 = MASTER_HREADY[5];

    end
    
  //===================================================================================================
  // MASTER 6
  //===================================================================================================
  if ( NUM_MASTERS > 6)
    begin  
      //output to master converter

      assign  MASTER_ARID[(6+1)*ID_WIDTH-1:6*ID_WIDTH]                                          = MASTER6_ARID;
      assign  MASTER_ARADDR[(6+1)*ADDR_WIDTH-1:6*ADDR_WIDTH]                                    = MASTER6_ARADDR;
      assign  MASTER_ARLEN[(6+1)*8-1:6*8]                                                       = MASTER6_ARLEN;
      assign  MASTER_ARSIZE[(6+1)*3-1:6*3]                                                      = MASTER6_ARSIZE;
      assign  MASTER_ARBURST[(6+1)*2-1:6*2]                                                     = MASTER6_ARBURST;
      assign  MASTER_ARLOCK[(6+1)*2-1:6*2]                                                      = MASTER6_ARLOCK;
      assign  MASTER_ARCACHE[(6+1)*4-1:6*4]                                                     = MASTER6_ARCACHE;
      assign  MASTER_ARPROT[(6+1)*3-1:6*3]                                                      = MASTER6_ARPROT;
      assign  MASTER_ARREGION[(6+1)*4-1:6*4]                                                    = MOD_MASTER6_ARREGION;
      assign  MASTER_ARQOS[(6+1)*4-1:6*4]                                                       = MOD_MASTER6_ARQOS;
      assign  MASTER_ARUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH]                                    = MASTER6_ARUSER;
      assign  MASTER_ARVALID[6]                                                                 = MASTER6_ARVALID;
      assign  MASTER_AWQOS[(6+1)*4-1:6*4]                                                       = MOD_MASTER6_AWQOS;
      assign  MASTER_AWREGION[(6+1)*4-1:6*4]                                                    = MOD_MASTER6_AWREGION;
      assign  MASTER_AWID[(6+1)*ID_WIDTH-1:6*ID_WIDTH]                                          = MASTER6_AWID;  
      assign  MASTER_AWADDR[(6+1)*ADDR_WIDTH-1:6*ADDR_WIDTH]                                    = MASTER6_AWADDR;  
      assign  MASTER_AWLEN[(6+1)*8-1:6*8]                                                       = MASTER6_AWLEN;  
      assign  MASTER_AWSIZE[(6+1)*3-1:6*3]                                                      = MASTER6_AWSIZE;  
      assign  MASTER_AWBURST[(6+1)*2-1:6*2]                                                     = MASTER6_AWBURST;  
      assign  MASTER_AWLOCK[(6+1)*2-1:6*2]                                                      = MASTER6_AWLOCK;  
      assign  MASTER_AWCACHE[(6+1)*4-1:6*4]                                                     = MASTER6_AWCACHE;  
      assign  MASTER_AWPROT[(6+1)*3-1:6*3]                                                      = MASTER6_AWPROT;  
      assign  MASTER_AWUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH]                                    = MASTER6_AWUSER;  
      assign  MASTER_AWVALID[6]                                                                 = MASTER6_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(6+1)*13-1:13*6]-1:MDW_LOWER_VEC[(6+1)*13-1:13*6]]     = MASTER6_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(6+1)*13-1:13*6]/8-1:MDW_LOWER_VEC[(6+1)*13-1:13*6]/8] = MASTER6_WSTRB;  
      assign  MASTER_WLAST[6]                                                                   = MASTER6_WLAST;  
      assign  MASTER_WUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH]                                     = MASTER6_WUSER;  
      assign  MASTER_WVALID[6]                                                                  = MASTER6_WVALID;  
      assign  MASTER_BREADY[6]                                                                  = MASTER6_BREADY;  
      assign  MASTER_RREADY[6]                                                                  = MASTER6_RREADY;

      assign MASTER6_RID        = MASTER_RID[(6+1)*ID_WIDTH-1:6*ID_WIDTH];
      assign MASTER6_RDATA      = MASTER_RDATA[MDW_UPPER_VEC[(6+1)*13-1:13*6]-1:MDW_LOWER_VEC[(6+1)*13-1:13*6]];
      assign MASTER6_RRESP      = MASTER_RRESP[(6+1)*2-1:6*2];
      assign MASTER6_RUSER      = MASTER_RUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH];
      assign MASTER6_BID        = MASTER_BID[(6+1)*ID_WIDTH-1:6*ID_WIDTH];
      assign MASTER6_BRESP      = MASTER_BRESP[(6+1)*2-1:6*2];
      assign MASTER6_BUSER      = MASTER_BUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH];
      assign MASTER6_ARREADY    = MASTER_ARREADY[6];
      assign MASTER6_RLAST      = MASTER_RLAST[6];
      assign MASTER6_RVALID     = MASTER_RVALID[6];
      assign MASTER6_AWREADY    = MASTER_AWREADY[6];
      assign MASTER6_WREADY     = MASTER_WREADY[6];
      assign MASTER6_BVALID     = MASTER_BVALID[6];

      // AHB interface
      assign MASTER_HADDR[32*(6+1)-1:32*6]                                                  = MASTER6_HADDR;
      assign MASTER_HBURST[3*(6+1)-1:3*6]                                                   = MASTER6_HBURST;
      assign MASTER_HMASTLOCK[6]                                                            = MASTER6_HMASTLOCK;
      assign MASTER_HPROT[7*(6+1)-1:7*6]                                                    = MASTER6_HPROT;          
      assign MASTER_HSIZE[3*(6+1)-1:3*6]                                                    = MASTER6_HSIZE;
      assign MASTER_HNONSEC[6]                                                              = MASTER6_HNONSEC;
      assign MASTER_HTRANS[2*(6+1)-1:2*6]                                                   = MASTER6_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(6+1)*13-1:13*6]-1:MDW_LOWER_VEC[(6+1)*13-1:13*6]] = MASTER6_HWDATA;
      assign MASTER6_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(6+1)*13-1:13*6]-1:MDW_LOWER_VEC[(6+1)*13-1:13*6]];
      assign MASTER_HWRITE[6]                                                               = MASTER6_HWRITE;
      assign MASTER6_HRESP                                                                  = MASTER_HRESP[6];
//      assign MASTER6_HEXOKAY                                                              = MASTER_HEXOKAY[6];
//      assign MASTER_HEXCL[6]                                                              = MASTER6_HEXCL;
      assign MASTER_HSEL[6]                                                                 = MASTER6_HSEL;
      assign MASTER6_HREADY                                                                 = MASTER_HREADY[6];

    end
    
  //===================================================================================================
  // MASTER 7
  //===================================================================================================
  if ( NUM_MASTERS > 7 )
    begin  
      //output to master converter
      
      assign  MASTER_ARID[(7+1)*ID_WIDTH-1:7*ID_WIDTH]                                          = MASTER7_ARID;
      assign  MASTER_ARADDR[(7+1)*ADDR_WIDTH-1:7*ADDR_WIDTH]                                    = MASTER7_ARADDR;
      assign  MASTER_ARLEN[(7+1)*8-1:7*8]                                                       = MASTER7_ARLEN;
      assign  MASTER_ARSIZE[(7+1)*3-1:7*3]                                                      = MASTER7_ARSIZE;
      assign  MASTER_ARBURST[(7+1)*2-1:7*2]                                                     = MASTER7_ARBURST;
      assign  MASTER_ARLOCK[(7+1)*2-1:7*2]                                                      = MASTER7_ARLOCK;
      assign  MASTER_ARCACHE[(7+1)*4-1:7*4]                                                     = MASTER7_ARCACHE;
      assign  MASTER_ARPROT[(7+1)*3-1:7*3]                                                      = MASTER7_ARPROT;
      assign  MASTER_ARREGION[(7+1)*4-1:7*4]                                                    = MOD_MASTER7_ARREGION;
      assign  MASTER_ARQOS[(7+1)*4-1:7*4]                                                       = MOD_MASTER7_ARQOS;
      assign  MASTER_ARUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH]                                    = MASTER7_ARUSER;
      assign  MASTER_ARVALID[7]                                                                 = MASTER7_ARVALID;
      assign  MASTER_AWQOS[(7+1)*4-1:7*4]                                                       = MOD_MASTER7_AWQOS;
      assign  MASTER_AWREGION[(7+1)*4-1:7*4]                                                    = MOD_MASTER7_AWREGION;
      assign  MASTER_AWID[(7+1)*ID_WIDTH-1:7*ID_WIDTH]                                          = MASTER7_AWID;  
      assign  MASTER_AWADDR[(7+1)*ADDR_WIDTH-1:7*ADDR_WIDTH]                                    = MASTER7_AWADDR;  
      assign  MASTER_AWLEN[(7+1)*8-1:7*8]                                                       = MASTER7_AWLEN;  
      assign  MASTER_AWSIZE[(7+1)*3-1:7*3]                                                      = MASTER7_AWSIZE;  
      assign  MASTER_AWBURST[(7+1)*2-1:7*2]                                                     = MASTER7_AWBURST;  
      assign  MASTER_AWLOCK[(7+1)*2-1:7*2]                                                      = MASTER7_AWLOCK;  
      assign  MASTER_AWCACHE[(7+1)*4-1:7*4]                                                     = MASTER7_AWCACHE;  
      assign  MASTER_AWPROT[(7+1)*3-1:7*3]                                                      = MASTER7_AWPROT;  
      assign  MASTER_AWUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH]                                    = MASTER7_AWUSER;  
      assign  MASTER_AWVALID[7]                                                                 = MASTER7_AWVALID;  
      assign  MASTER_WDATA[MDW_UPPER_VEC[(7+1)*13-1:13*7]-1:MDW_LOWER_VEC[(7+1)*13-1:13*7]]     = MASTER7_WDATA;  
      assign  MASTER_WSTRB[MDW_UPPER_VEC[(7+1)*13-1:13*7]/8-1:MDW_LOWER_VEC[(7+1)*13-1:13*7]/8] = MASTER7_WSTRB;  
      assign  MASTER_WLAST[7]                                                                   = MASTER7_WLAST;  
      assign  MASTER_WUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH]                                     = MASTER7_WUSER;  
      assign  MASTER_WVALID[7]                                                                  = MASTER7_WVALID;  
      assign  MASTER_BREADY[7]                                                                  = MASTER7_BREADY;  
      assign  MASTER_RREADY[7]                                                                  = MASTER7_RREADY;

      assign   MASTER7_RID      = MASTER_RID[(7+1)*ID_WIDTH-1:7*ID_WIDTH];
      assign   MASTER7_RDATA    = MASTER_RDATA[MDW_UPPER_VEC[(7+1)*13-1:13*7]-1:MDW_LOWER_VEC[(7+1)*13-1:13*7]];
      assign   MASTER7_RRESP    = MASTER_RRESP[(7+1)*2-1:7*2];
      assign   MASTER7_RUSER    = MASTER_RUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH];
      assign   MASTER7_BID      = MASTER_BID[(7+1)*ID_WIDTH-1:7*ID_WIDTH];
      assign   MASTER7_BRESP    = MASTER_BRESP[(7+1)*2-1:7*2];
      assign   MASTER7_BUSER    = MASTER_BUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH];
      assign   MASTER7_ARREADY  = MASTER_ARREADY[7];
      assign   MASTER7_RLAST    = MASTER_RLAST[7];
      assign   MASTER7_RVALID   = MASTER_RVALID[7];
      assign   MASTER7_AWREADY  = MASTER_AWREADY[7];
      assign   MASTER7_WREADY   = MASTER_WREADY[7];
      assign   MASTER7_BVALID   = MASTER_BVALID[7];

      // AHB interface
      assign MASTER_HADDR[32*(7+1)-1:32*7]                                                  = MASTER7_HADDR;
      assign MASTER_HBURST[3*(7+1)-1:3*7]                                                   = MASTER7_HBURST;
      assign MASTER_HMASTLOCK[7]                                                            = MASTER7_HMASTLOCK;
      assign MASTER_HPROT[7*(7+1)-1:7*7]                                                    = MASTER7_HPROT;          
      assign MASTER_HSIZE[3*(7+1)-1:3*7]                                                    = MASTER7_HSIZE;
      assign MASTER_HNONSEC[7]                                                              = MASTER7_HNONSEC;
      assign MASTER_HTRANS[2*(7+1)-1:2*7]                                                   = MASTER7_HTRANS;
      assign MASTER_HWDATA[MDW_UPPER_VEC[(7+1)*13-1:13*7]-1:MDW_LOWER_VEC[(7+1)*13-1:13*7]] = MASTER7_HWDATA;
      assign MASTER7_HRDATA                                                                 = MASTER_HRDATA[MDW_UPPER_VEC[(7+1)*13-1:13*7]-1:MDW_LOWER_VEC[(7+1)*13-1:13*7]];
      assign MASTER_HWRITE[7]                                                               = MASTER7_HWRITE;
      assign MASTER7_HRESP                                                                  = MASTER_HRESP[7];
//      assign MASTER7_HEXOKAY                                                              = MASTER_HEXOKAY[7];
//      assign MASTER_HEXCL[7]                                                              = MASTER7_HEXCL;
      assign MASTER_HSEL[7]                                                                 = MASTER7_HSEL;
      assign MASTER7_HREADY                                                                 = MASTER_HREADY[7];

    end
      
  //===================================================================
  //Slave0 Combine Signals
  //===================================================================
  //======================= SLAVE0 TO/FROM External Side=================
  //Outputs
  //
  assign  SLAVE0_AWID     = SLAVE_AWID[(0+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
  assign  SLAVE0_AWADDR   = SLAVE_AWADDR[(0+1)*ADDR_WIDTH-1:0*ADDR_WIDTH];  
  assign  SLAVE0_AWLEN    = SLAVE_AWLEN[(0+1)*8-1:0*8];  
  assign  SLAVE0_AWSIZE   = SLAVE_AWSIZE[(0+1)*3-1:0*3];  
  assign  SLAVE0_AWBURST  = SLAVE_AWBURST[(0+1)*2-1:0*2];  
  assign  SLAVE0_AWLOCK   = SLAVE_AWLOCK[(0+1)*2-1:0*2];  
  assign  SLAVE0_AWCACHE  = SLAVE_AWCACHE[(0+1)*4-1:0*4];  
  assign  SLAVE0_AWPROT   = SLAVE_AWPROT[(0+1)*3-1:0*3];  
  assign  SLAVE0_AWREGION = SLAVE_AWREGION[(0+1)*4-1:0*4];   
  assign  SLAVE0_AWQOS    = SLAVE_AWQOS[(0+1)*4-1:0*4];  
  assign  SLAVE0_AWUSER   = SLAVE_AWUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH];  
  assign  SLAVE0_AWVALID  = SLAVE_AWVALID[0];  
  assign  SLAVE0_WID      = SLAVE_WID[(0+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
  assign  SLAVE0_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(0+1)*13-1:13*0]-1:SDW_LOWER_VEC[(0+1)*13-1:13*0]];  
  assign  SLAVE0_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(0+1)*13-1:13*0]/8-1:SDW_LOWER_VEC[(0+1)*13-1:13*0]];  
  assign  SLAVE0_WLAST    = SLAVE_WLAST[0];  
  assign  SLAVE0_WUSER    = SLAVE_WUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH];  
  assign  SLAVE0_WVALID   = SLAVE_WVALID[0];      
  assign  SLAVE0_BREADY   = SLAVE_BREADY[0];        
  assign  SLAVE0_ARID     = SLAVE_ARID[(0+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
  assign  SLAVE0_ARADDR   = SLAVE_ARADDR[(0+1)*ADDR_WIDTH-1:0*ADDR_WIDTH];  
  assign  SLAVE0_ARLEN    = SLAVE_ARLEN[(0+1)*8-1:0*8];  
  assign  SLAVE0_ARSIZE   = SLAVE_ARSIZE[(0+1)*3-1:0*3];  
  assign  SLAVE0_ARBURST  = SLAVE_ARBURST[(0+1)*2-1:0*2];  
  assign  SLAVE0_ARLOCK   = SLAVE_ARLOCK[(0+1)*2-1:0*2];  
  assign  SLAVE0_ARCACHE  = SLAVE_ARCACHE[(0+1)*4-1:0*4] ;  
  assign  SLAVE0_ARPROT   = SLAVE_ARPROT[(0+1)*3-1:0*3] ;  
  assign  SLAVE0_ARREGION = SLAVE_ARREGION[(0+1)*4-1:0*4];   
  assign  SLAVE0_ARQOS    = SLAVE_ARQOS[(0+1)*4-1:0*4];  
  assign  SLAVE0_ARUSER   = SLAVE_ARUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH];  
  assign  SLAVE0_ARVALID  = SLAVE_ARVALID[0];      
  assign  SLAVE0_RREADY   = SLAVE_RREADY[0];  

  //Inputs      
  assign  SLAVE_AWREADY[0]                                                                 = SLAVE0_AWREADY;          
  assign  SLAVE_WREADY[0]                                                                  = SLAVE0_WREADY;        
  assign  SLAVE_BID[(0+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE0_BID;  
  assign  SLAVE_BRESP[(0+1)*2-1:0*2]                                                       = SLAVE0_BRESP;  
  assign  SLAVE_BUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH]                                     = SLAVE0_BUSER;  
  assign  SLAVE_BVALID[0]                                                                  = SLAVE0_BVALID;        
  assign  SLAVE_ARREADY[0]                                                                 = SLAVE0_ARREADY;        
  assign  SLAVE_RID[(0+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:0*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE0_RID;  
  assign  SLAVE_RDATA[SDW_UPPER_VEC[(0+1)*13-1:13*0]-1:SDW_LOWER_VEC[(0+1)*13-1:13*0]]     = SLAVE0_RDATA;  
  assign  SLAVE_RRESP[(0+1)*2-1:0*2]                                                       = SLAVE0_RRESP;  
  assign  SLAVE_RLAST[0]                                                                   = SLAVE0_RLAST;  
  assign  SLAVE_RUSER[(0+1)*USER_WIDTH-1:0*USER_WIDTH]                                     = SLAVE0_RUSER;  
  assign  SLAVE_RVALID[0]                                                                  = SLAVE0_RVALID;

  if ( NUM_SLAVES > 1 )
    begin
      //===================================================================
      //Slave1 Combine Signals
      //===================================================================
      //======================= SLAVE1 TO/FROM External Side=================
      //Outputs
      //
      assign  SLAVE1_AWID     = SLAVE_AWID[(1+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:1*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE1_AWADDR   = SLAVE_AWADDR[(1+1)*ADDR_WIDTH-1:1*ADDR_WIDTH];  
      assign  SLAVE1_AWLEN    = SLAVE_AWLEN[(1+1)*8-1:1*8];  
      assign  SLAVE1_AWSIZE   = SLAVE_AWSIZE[(1+1)*3-1:1*3];  
      assign  SLAVE1_AWBURST  = SLAVE_AWBURST[(1+1)*2-1:1*2];  
      assign  SLAVE1_AWLOCK   = SLAVE_AWLOCK[(1+1)*2-1:1*2];  
      assign  SLAVE1_AWCACHE  = SLAVE_AWCACHE[(1+1)*4-1:1*4];  
      assign  SLAVE1_AWPROT   = SLAVE_AWPROT[(1+1)*3-1:1*3];  
      assign  SLAVE1_AWREGION = SLAVE_AWREGION[(1+1)*4-1:1*4];   
      assign  SLAVE1_AWQOS    = SLAVE_AWQOS[(1+1)*4-1:1*4];  
      assign  SLAVE1_AWUSER   = SLAVE_AWUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH];  
      assign  SLAVE1_AWVALID  = SLAVE_AWVALID[1];        
      assign  SLAVE1_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(1+1)*13-1:13*1]-1:SDW_LOWER_VEC[(1+1)*13-1:13*1]];  
      assign  SLAVE1_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(1+1)*13-1:13*1]/8-1:SDW_LOWER_VEC[(1+1)*13-1:13*1]/8];  
      assign  SLAVE1_WLAST    = SLAVE_WLAST[1];  
      assign  SLAVE1_WID      = SLAVE_WID[(1+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:1*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE1_WUSER    = SLAVE_WUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH];  
      assign  SLAVE1_WVALID   = SLAVE_WVALID[1];      
      assign  SLAVE1_BREADY   = SLAVE_BREADY[1];        
      assign  SLAVE1_ARID     = SLAVE_ARID[(1+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:1*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE1_ARADDR   = SLAVE_ARADDR[(1+1)*ADDR_WIDTH-1:1*ADDR_WIDTH];  
      assign  SLAVE1_ARLEN    = SLAVE_ARLEN[(1+1)*8-1:1*8];  
      assign  SLAVE1_ARSIZE   = SLAVE_ARSIZE[(1+1)*3-1:1*3];  
      assign  SLAVE1_ARBURST  = SLAVE_ARBURST[(1+1)*2-1:1*2];  
      assign  SLAVE1_ARLOCK   = SLAVE_ARLOCK[(1+1)*2-1:1*2];  
      assign  SLAVE1_ARCACHE  = SLAVE_ARCACHE[(1+1)*4-1:1*4] ;  
      assign  SLAVE1_ARPROT   = SLAVE_ARPROT[(1+1)*3-1:1*3] ;  
      assign  SLAVE1_ARREGION = SLAVE_ARREGION[(1+1)*4-1:1*4];   
      assign  SLAVE1_ARQOS    = SLAVE_ARQOS[(1+1)*4-1:1*4];  
      assign  SLAVE1_ARUSER   = SLAVE_ARUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH];  
      assign  SLAVE1_ARVALID  = SLAVE_ARVALID[1];      
      assign  SLAVE1_RREADY   = SLAVE_RREADY[1];  

      //Inputs      
      assign  SLAVE_AWREADY[1]                                                                 = SLAVE1_AWREADY;          
      assign  SLAVE_WREADY[1]                                                                  = SLAVE1_WREADY;        
      assign  SLAVE_BID[(1+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:1*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE1_BID;  
      assign  SLAVE_BRESP[(1+1)*2-1:1*2]                                                       = SLAVE1_BRESP;  
      assign  SLAVE_BUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH]                                     = SLAVE1_BUSER;  
      assign  SLAVE_BVALID[1]                                                                  = SLAVE1_BVALID;        
      assign  SLAVE_ARREADY[1]                                                                 = SLAVE1_ARREADY;        
      assign  SLAVE_RID[(1+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:1*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE1_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(1+1)*13-1:13*1]-1:SDW_LOWER_VEC[(1+1)*13-1:13*1]]     = SLAVE1_RDATA;  
      assign  SLAVE_RRESP[(1+1)*2-1:1*2]                                                       = SLAVE1_RRESP;  
      assign  SLAVE_RLAST[1]                                                                   = SLAVE1_RLAST;  
      assign  SLAVE_RUSER[(1+1)*USER_WIDTH-1:1*USER_WIDTH]                                     = SLAVE1_RUSER;  
      assign  SLAVE_RVALID[1]                                                                  = SLAVE1_RVALID;
    end
    
  if ( NUM_SLAVES > 2 )
    begin
      //===================================================================
      //Slave2 Combine Signals
      //===================================================================
      //======================= SLAVE2 TO/FROM External Side=================
      //Outputs
      //
      assign  SLAVE2_AWID     = SLAVE_AWID[(2+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:2*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE2_AWADDR   = SLAVE_AWADDR[(2+1)*ADDR_WIDTH-1:2*ADDR_WIDTH];  
      assign  SLAVE2_AWLEN    = SLAVE_AWLEN[(2+1)*8-1:2*8];  
      assign  SLAVE2_AWSIZE   = SLAVE_AWSIZE[(2+1)*3-1:2*3];  
      assign  SLAVE2_AWBURST  = SLAVE_AWBURST[(2+1)*2-1:2*2];  
      assign  SLAVE2_AWLOCK   = SLAVE_AWLOCK[(2+1)*2-1:2*2];  
      assign  SLAVE2_AWCACHE  = SLAVE_AWCACHE[(2+1)*4-1:2*4];  
      assign  SLAVE2_AWPROT   = SLAVE_AWPROT[(2+1)*3-1:2*3];  
      assign  SLAVE2_AWREGION = SLAVE_AWREGION[(2+1)*4-1:2*4];   
      assign  SLAVE2_AWQOS    = SLAVE_AWQOS[(2+1)*4-1:2*4];  
      assign  SLAVE2_AWUSER   = SLAVE_AWUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH];  
      assign  SLAVE2_AWVALID  = SLAVE_AWVALID[2];
      assign  SLAVE2_WID      = SLAVE_WID[(2+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:2*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE2_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(2+1)*13-1:13*2]-1:SDW_LOWER_VEC[(2+1)*13-1:13*2]];  
      assign  SLAVE2_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(2+1)*13-1:13*2]/8-1:SDW_LOWER_VEC[(2+1)*13-1:13*2]/8];  
      assign  SLAVE2_WLAST    = SLAVE_WLAST[2];  
      assign  SLAVE2_WUSER    = SLAVE_WUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH];  
      assign  SLAVE2_WVALID   = SLAVE_WVALID[2];      
      assign  SLAVE2_BREADY   = SLAVE_BREADY[2];        
      assign  SLAVE2_ARID     = SLAVE_ARID[(2+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:2*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE2_ARADDR   = SLAVE_ARADDR[(2+1)*ADDR_WIDTH-1:2*ADDR_WIDTH];  
      assign  SLAVE2_ARLEN    = SLAVE_ARLEN[(2+1)*8-1:2*8];  
      assign  SLAVE2_ARSIZE   = SLAVE_ARSIZE[(2+1)*3-1:2*3];  
      assign  SLAVE2_ARBURST  = SLAVE_ARBURST[(2+1)*2-1:2*2];  
      assign  SLAVE2_ARLOCK   = SLAVE_ARLOCK[(2+1)*2-1:2*2];  
      assign  SLAVE2_ARCACHE  = SLAVE_ARCACHE[(2+1)*4-1:2*4] ;  
      assign  SLAVE2_ARPROT   = SLAVE_ARPROT[(2+1)*3-1:2*3] ;  
      assign  SLAVE2_ARREGION = SLAVE_ARREGION[(2+1)*4-1:2*4];   
      assign  SLAVE2_ARQOS    = SLAVE_ARQOS[(2+1)*4-1:2*4];  
      assign  SLAVE2_ARUSER   = SLAVE_ARUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH];  
      assign  SLAVE2_ARVALID  = SLAVE_ARVALID[2];      
      assign  SLAVE2_RREADY   = SLAVE_RREADY[2];  

      //Inputs      
      assign  SLAVE_AWREADY[2]                                                                 = SLAVE2_AWREADY;          
      assign  SLAVE_WREADY[2]                                                                  = SLAVE2_WREADY;        
      assign  SLAVE_BID[(2+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:2*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE2_BID;  
      assign  SLAVE_BRESP[(2+1)*2-1:2*2]                                                       = SLAVE2_BRESP;  
      assign  SLAVE_BUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH]                                     = SLAVE2_BUSER;  
      assign  SLAVE_BVALID[2]                                                                  = SLAVE2_BVALID;        
      assign  SLAVE_ARREADY[2]                                                                 = SLAVE2_ARREADY;        
      assign  SLAVE_RID[(2+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:2*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE2_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(2+1)*13-1:13*2]-1:SDW_LOWER_VEC[(2+1)*13-1:13*2]]     = SLAVE2_RDATA;  
      assign  SLAVE_RRESP[(2+1)*2-1:2*2]                                                       = SLAVE2_RRESP;  
      assign  SLAVE_RLAST[2]                                                                   = SLAVE2_RLAST;  
      assign  SLAVE_RUSER[(2+1)*USER_WIDTH-1:2*USER_WIDTH]                                     = SLAVE2_RUSER;  
      assign  SLAVE_RVALID[2]                                                                  = SLAVE2_RVALID;
    end
    
  if ( NUM_SLAVES > 3 )
    begin    
      //===================================================================
      //Slave3 Combine Signals
      //===================================================================
      //======================= SLAVE3 TO/FROM External Side=================
      //Outputs
      assign  SLAVE3_AWID     = SLAVE_AWID[(3+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:3*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE3_AWADDR   = SLAVE_AWADDR[(3+1)*ADDR_WIDTH-1:3*ADDR_WIDTH];  
      assign  SLAVE3_AWLEN    = SLAVE_AWLEN[(3+1)*8-1:3*8];  
      assign  SLAVE3_AWSIZE   = SLAVE_AWSIZE[(3+1)*3-1:3*3];  
      assign  SLAVE3_AWBURST  = SLAVE_AWBURST[(3+1)*2-1:3*2];  
      assign  SLAVE3_AWLOCK   = SLAVE_AWLOCK[(3+1)*2-1:3*2];  
      assign  SLAVE3_AWCACHE  = SLAVE_AWCACHE[(3+1)*4-1:3*4];  
      assign  SLAVE3_AWPROT   = SLAVE_AWPROT[(3+1)*3-1:3*3];  
      assign  SLAVE3_AWREGION = SLAVE_AWREGION[(3+1)*4-1:3*4];   
      assign  SLAVE3_AWQOS    = SLAVE_AWQOS[(3+1)*4-1:3*4];  
      assign  SLAVE3_AWUSER   = SLAVE_AWUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH];  
      assign  SLAVE3_AWVALID  = SLAVE_AWVALID[3];        
      assign  SLAVE3_WID      = SLAVE_WID[(3+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:3*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE3_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(3+1)*13-1:13*3]-1:SDW_LOWER_VEC[(3+1)*13-1:13*3]];  
      assign  SLAVE3_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(3+1)*13-1:13*3]/8-1:SDW_LOWER_VEC[(3+1)*13-1:13*3]/8];  
      assign  SLAVE3_WLAST    = SLAVE_WLAST[3];  
      assign  SLAVE3_WUSER    = SLAVE_WUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH];  
      assign  SLAVE3_WVALID   = SLAVE_WVALID[3];      
      assign  SLAVE3_BREADY   = SLAVE_BREADY[3];        
      assign  SLAVE3_ARID     = SLAVE_ARID[(3+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:3*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE3_ARADDR   = SLAVE_ARADDR[(3+1)*ADDR_WIDTH-1:3*ADDR_WIDTH];  
      assign  SLAVE3_ARLEN    = SLAVE_ARLEN[(3+1)*8-1:3*8];  
      assign  SLAVE3_ARSIZE   = SLAVE_ARSIZE[(3+1)*3-1:3*3];  
      assign  SLAVE3_ARBURST  = SLAVE_ARBURST[(3+1)*2-1:3*2];  
      assign  SLAVE3_ARLOCK   = SLAVE_ARLOCK[(3+1)*2-1:3*2];  
      assign  SLAVE3_ARCACHE  = SLAVE_ARCACHE[(3+1)*4-1:3*4] ;  
      assign  SLAVE3_ARPROT   = SLAVE_ARPROT[(3+1)*3-1:3*3] ;  
      assign  SLAVE3_ARREGION = SLAVE_ARREGION[(3+1)*4-1:3*4];   
      assign  SLAVE3_ARQOS    = SLAVE_ARQOS[(3+1)*4-1:3*4];  
      assign  SLAVE3_ARUSER   = SLAVE_ARUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH];  
      assign  SLAVE3_ARVALID  = SLAVE_ARVALID[3];      
      assign  SLAVE3_RREADY   = SLAVE_RREADY[3];  

      //Inputs      
      assign  SLAVE_AWREADY[3]                                                                 = SLAVE3_AWREADY;          
      assign  SLAVE_WREADY[3]                                                                  = SLAVE3_WREADY;        
      assign  SLAVE_BID[(3+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:3*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE3_BID;  
      assign  SLAVE_BRESP[(3+1)*2-1:3*2]                                                       = SLAVE3_BRESP;  
      assign  SLAVE_BUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH]                                     = SLAVE3_BUSER;  
      assign  SLAVE_BVALID[3]                                                                  = SLAVE3_BVALID;        
      assign  SLAVE_ARREADY[3]                                                                 = SLAVE3_ARREADY;        
      assign  SLAVE_RID[(3+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:3*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE3_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(3+1)*13-1:13*3]-1:SDW_LOWER_VEC[(3+1)*13-1:13*3]]     = SLAVE3_RDATA;  
      assign  SLAVE_RRESP[(3+1)*2-1:3*2]                                                       = SLAVE3_RRESP;  
      assign  SLAVE_RLAST[3]                                                                   = SLAVE3_RLAST;  
      assign  SLAVE_RUSER[(3+1)*USER_WIDTH-1:3*USER_WIDTH]                                     = SLAVE3_RUSER;  
      assign  SLAVE_RVALID[3]                                                                  = SLAVE3_RVALID;
    end
    
  if ( NUM_SLAVES > 4 )
    begin
      //===================================================================
      //Slave4 Combine Signals
      //===================================================================
      //======================= SLAVE4 TO/FROM External Side=================
      //Outputs
      //
      assign  SLAVE4_AWID     = SLAVE_AWID[(4+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:4*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE4_AWADDR   = SLAVE_AWADDR[(4+1)*ADDR_WIDTH-1:4*ADDR_WIDTH];  
      assign  SLAVE4_AWLEN    = SLAVE_AWLEN[(4+1)*8-1:4*8];  
      assign  SLAVE4_AWSIZE   = SLAVE_AWSIZE[(4+1)*3-1:4*3];  
      assign  SLAVE4_AWBURST  = SLAVE_AWBURST[(4+1)*2-1:4*2];  
      assign  SLAVE4_AWLOCK   = SLAVE_AWLOCK[(4+1)*2-1:4*2];  
      assign  SLAVE4_AWCACHE  = SLAVE_AWCACHE[(4+1)*4-1:4*4];  
      assign  SLAVE4_AWPROT   = SLAVE_AWPROT[(4+1)*3-1:4*3];  
      assign  SLAVE4_AWREGION = SLAVE_AWREGION[(4+1)*4-1:4*4];   
      assign  SLAVE4_AWQOS    = SLAVE_AWQOS[(4+1)*4-1:4*4];  
      assign  SLAVE4_AWUSER   = SLAVE_AWUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH];  
      assign  SLAVE4_AWVALID  = SLAVE_AWVALID[4];  
      assign  SLAVE4_WID      = SLAVE_WID[(4+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:4*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE4_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(4+1)*13-1:13*4]-1:SDW_LOWER_VEC[(4+1)*13-1:13*4]];  
      assign  SLAVE4_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(4+1)*13-1:13*4]/8-1:SDW_LOWER_VEC[(4+1)*13-1:13*4]/8];  
      assign  SLAVE4_WLAST    = SLAVE_WLAST[4];  
      assign  SLAVE4_WUSER    = SLAVE_WUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH];  
      assign  SLAVE4_WVALID   = SLAVE_WVALID[4];      
      assign  SLAVE4_BREADY   = SLAVE_BREADY[4];        
      assign  SLAVE4_ARID     = SLAVE_ARID[(4+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:4*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE4_ARADDR   = SLAVE_ARADDR[(4+1)*ADDR_WIDTH-1:4*ADDR_WIDTH];  
      assign  SLAVE4_ARLEN    = SLAVE_ARLEN[(4+1)*8-1:4*8];  
      assign  SLAVE4_ARSIZE   = SLAVE_ARSIZE[(4+1)*3-1:4*3];  
      assign  SLAVE4_ARBURST  = SLAVE_ARBURST[(4+1)*2-1:4*2];  
      assign  SLAVE4_ARLOCK   = SLAVE_ARLOCK[(4+1)*2-1:4*2];  
      assign  SLAVE4_ARCACHE  = SLAVE_ARCACHE[(4+1)*4-1:4*4] ;  
      assign  SLAVE4_ARPROT   = SLAVE_ARPROT[(4+1)*3-1:4*3] ;  
      assign  SLAVE4_ARREGION = SLAVE_ARREGION[(4+1)*4-1:4*4];   
      assign  SLAVE4_ARQOS    = SLAVE_ARQOS[(4+1)*4-1:4*4];  
      assign  SLAVE4_ARUSER   = SLAVE_ARUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH];  
      assign  SLAVE4_ARVALID  = SLAVE_ARVALID[4];      
      assign  SLAVE4_RREADY   = SLAVE_RREADY[4];  

      //Inputs      
      assign  SLAVE_AWREADY[4]                                                                 = SLAVE4_AWREADY;          
      assign  SLAVE_WREADY[4]                                                                  = SLAVE4_WREADY;        
      assign  SLAVE_BID[(4+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:4*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE4_BID;  
      assign  SLAVE_BRESP[(4+1)*2-1:4*2]                                                       = SLAVE4_BRESP;  
      assign  SLAVE_BUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH]                                     = SLAVE4_BUSER;  
      assign  SLAVE_BVALID[4]                                                                  = SLAVE4_BVALID;        
      assign  SLAVE_ARREADY[4]                                                                 = SLAVE4_ARREADY;        
      assign  SLAVE_RID[(4+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:4*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE4_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(4+1)*13-1:13*4]-1:SDW_LOWER_VEC[(4+1)*13-1:13*4]]     = SLAVE4_RDATA;  
      assign  SLAVE_RRESP[(4+1)*2-1:4*2]                                                       = SLAVE4_RRESP;  
      assign  SLAVE_RLAST[4]                                                                   = SLAVE4_RLAST;  
      assign  SLAVE_RUSER[(4+1)*USER_WIDTH-1:4*USER_WIDTH]                                     = SLAVE4_RUSER;  
      assign  SLAVE_RVALID[4]                                                                  = SLAVE4_RVALID;
    end
    
  if ( NUM_SLAVES > 5 )
    begin        
      //===================================================================
      //Slave5 Combine Signals
      //===================================================================
      //======================= SLAVE5 TO/FROM External Side=================
      //Outputs  
      assign  SLAVE5_AWID     = SLAVE_AWID[(5+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:5*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE5_AWADDR   = SLAVE_AWADDR[(5+1)*ADDR_WIDTH-1:5*ADDR_WIDTH];  
      assign  SLAVE5_AWLEN    = SLAVE_AWLEN[(5+1)*8-1:5*8];  
      assign  SLAVE5_AWSIZE   = SLAVE_AWSIZE[(5+1)*3-1:5*3];  
      assign  SLAVE5_AWBURST  = SLAVE_AWBURST[(5+1)*2-1:5*2];  
      assign  SLAVE5_AWLOCK   = SLAVE_AWLOCK[(5+1)*2-1:5*2];  
      assign  SLAVE5_AWCACHE  = SLAVE_AWCACHE[(5+1)*4-1:5*4];  
      assign  SLAVE5_AWPROT   = SLAVE_AWPROT[(5+1)*3-1:5*3];  
      assign  SLAVE5_AWREGION = SLAVE_AWREGION[(5+1)*4-1:5*4];   
      assign  SLAVE5_AWQOS    = SLAVE_AWQOS[(5+1)*4-1:5*4];  
      assign  SLAVE5_AWUSER   = SLAVE_AWUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH];  
      assign  SLAVE5_AWVALID  = SLAVE_AWVALID[5];
      assign  SLAVE5_WID      = SLAVE_WID[(5+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:5*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE5_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(5+1)*13-1:13*5]-1:SDW_LOWER_VEC[(5+1)*13-1:13*5]];  
      assign  SLAVE5_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(5+1)*13-1:13*5]/8-1:SDW_LOWER_VEC[(5+1)*13-1:13*5]/8];  
      assign  SLAVE5_WLAST    = SLAVE_WLAST[5];  
      assign  SLAVE5_WUSER    = SLAVE_WUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH];  
      assign  SLAVE5_WVALID   = SLAVE_WVALID[5];      
      assign  SLAVE5_BREADY   = SLAVE_BREADY[5];        
      assign  SLAVE5_ARID     = SLAVE_ARID[(5+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:5*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE5_ARADDR   = SLAVE_ARADDR[(5+1)*ADDR_WIDTH-1:5*ADDR_WIDTH];  
      assign  SLAVE5_ARLEN    = SLAVE_ARLEN[(5+1)*8-1:5*8];  
      assign  SLAVE5_ARSIZE   = SLAVE_ARSIZE[(5+1)*3-1:5*3];  
      assign  SLAVE5_ARBURST  = SLAVE_ARBURST[(5+1)*2-1:5*2];  
      assign  SLAVE5_ARLOCK   = SLAVE_ARLOCK[(5+1)*2-1:5*2];  
      assign  SLAVE5_ARCACHE  = SLAVE_ARCACHE[(5+1)*4-1:5*4] ;  
      assign  SLAVE5_ARPROT   = SLAVE_ARPROT[(5+1)*3-1:5*3] ;  
      assign  SLAVE5_ARREGION = SLAVE_ARREGION[(5+1)*4-1:5*4];   
      assign  SLAVE5_ARQOS    = SLAVE_ARQOS[(5+1)*4-1:5*4];  
      assign  SLAVE5_ARUSER   = SLAVE_ARUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH];  
      assign  SLAVE5_ARVALID  = SLAVE_ARVALID[5];      
      assign  SLAVE5_RREADY   = SLAVE_RREADY[5];  

      //Inputs      
      assign  SLAVE_AWREADY[5]                                                                 = SLAVE5_AWREADY;          
      assign  SLAVE_WREADY[5]                                                                  = SLAVE5_WREADY;        
      assign  SLAVE_BID[(5+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:5*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE5_BID;  
      assign  SLAVE_BRESP[(5+1)*2-1:5*2]                                                       = SLAVE5_BRESP;  
      assign  SLAVE_BUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH]                                     = SLAVE5_BUSER;  
      assign  SLAVE_BVALID[5]                                                                  = SLAVE5_BVALID;        
      assign  SLAVE_ARREADY[5]                                                                 = SLAVE5_ARREADY;        
      assign  SLAVE_RID[(5+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:5*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE5_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(5+1)*13-1:13*5]-1:SDW_LOWER_VEC[(5+1)*13-1:13*5]]     = SLAVE5_RDATA;  
      assign  SLAVE_RRESP[(5+1)*2-1:5*2]                                                       = SLAVE5_RRESP;  
      assign  SLAVE_RLAST[5]                                                                   = SLAVE5_RLAST;  
      assign  SLAVE_RUSER[(5+1)*USER_WIDTH-1:5*USER_WIDTH]                                     = SLAVE5_RUSER;  
      assign  SLAVE_RVALID[5]                                                                  = SLAVE5_RVALID;
    end
    
  if ( NUM_SLAVES > 6 )
    begin
      
      //===================================================================
      //Slave6 Combine Signals
      //===================================================================
      //======================= SLAVE6 TO/FROM External Side=================
      //Outputs
      assign  SLAVE6_AWID     = SLAVE_AWID[(6+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:6*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE6_AWADDR   = SLAVE_AWADDR[(6+1)*ADDR_WIDTH-1:6*ADDR_WIDTH];  
      assign  SLAVE6_AWLEN    = SLAVE_AWLEN[(6+1)*8-1:6*8];  
      assign  SLAVE6_AWSIZE   = SLAVE_AWSIZE[(6+1)*3-1:6*3];  
      assign  SLAVE6_AWBURST  = SLAVE_AWBURST[(6+1)*2-1:6*2];  
      assign  SLAVE6_AWLOCK   = SLAVE_AWLOCK[(6+1)*2-1:6*2];  
      assign  SLAVE6_AWCACHE  = SLAVE_AWCACHE[(6+1)*4-1:6*4];  
      assign  SLAVE6_AWPROT   = SLAVE_AWPROT[(6+1)*3-1:6*3];  
      assign  SLAVE6_AWREGION = SLAVE_AWREGION[(6+1)*4-1:6*4];   
      assign  SLAVE6_AWQOS    = SLAVE_AWQOS[(6+1)*4-1:6*4];  
      assign  SLAVE6_AWUSER   = SLAVE_AWUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH];  
      assign  SLAVE6_AWVALID  = SLAVE_AWVALID[6];  
      assign  SLAVE6_WID      = SLAVE_WID[(6+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:6*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE6_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(6+1)*13-1:13*6]-1:SDW_LOWER_VEC[(6+1)*13-1:13*6]];  
      assign  SLAVE6_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(6+1)*13-1:13*6]/8-1:SDW_LOWER_VEC[(6+1)*13-1:13*6]/8];  
      assign  SLAVE6_WLAST    = SLAVE_WLAST[6];  
      assign  SLAVE6_WUSER    = SLAVE_WUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH];  
      assign  SLAVE6_WVALID   = SLAVE_WVALID[6];      
      assign  SLAVE6_BREADY   = SLAVE_BREADY[6];        
      assign  SLAVE6_ARID     = SLAVE_ARID[(6+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:6*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE6_ARADDR   = SLAVE_ARADDR[(6+1)*ADDR_WIDTH-1:6*ADDR_WIDTH];  
      assign  SLAVE6_ARLEN    = SLAVE_ARLEN[(6+1)*8-1:6*8];  
      assign  SLAVE6_ARSIZE   = SLAVE_ARSIZE[(6+1)*3-1:6*3];  
      assign  SLAVE6_ARBURST  = SLAVE_ARBURST[(6+1)*2-1:6*2];  
      assign  SLAVE6_ARLOCK   = SLAVE_ARLOCK[(6+1)*2-1:6*2];  
      assign  SLAVE6_ARCACHE  = SLAVE_ARCACHE[(6+1)*4-1:6*4] ;  
      assign  SLAVE6_ARPROT   = SLAVE_ARPROT[(6+1)*3-1:6*3] ;  
      assign  SLAVE6_ARREGION = SLAVE_ARREGION[(6+1)*4-1:6*4];   
      assign  SLAVE6_ARQOS    = SLAVE_ARQOS[(6+1)*4-1:6*4];  
      assign  SLAVE6_ARUSER   = SLAVE_ARUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH];  
      assign  SLAVE6_ARVALID  = SLAVE_ARVALID[6];      
      assign  SLAVE6_RREADY   = SLAVE_RREADY[6];  

      //Inputs      
      assign  SLAVE_AWREADY[6]                                                                 = SLAVE6_AWREADY;          
      assign  SLAVE_WREADY[6]                                                                  = SLAVE6_WREADY;        
      assign  SLAVE_BID[(6+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:6*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE6_BID;  
      assign  SLAVE_BRESP[(6+1)*2-1:6*2]                                                       = SLAVE6_BRESP;  
      assign  SLAVE_BUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH]                                     = SLAVE6_BUSER;  
      assign  SLAVE_BVALID[6]                                                                  = SLAVE6_BVALID;        
      assign  SLAVE_ARREADY[6]                                                                 = SLAVE6_ARREADY;        
      assign  SLAVE_RID[(6+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:6*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE6_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(6+1)*13-1:13*6]-1:SDW_LOWER_VEC[(6+1)*13-1:13*6]]     = SLAVE6_RDATA;  
      assign  SLAVE_RRESP[(6+1)*2-1:6*2]                                                       = SLAVE6_RRESP;  
      assign  SLAVE_RLAST[6]                                                                   = SLAVE6_RLAST;  
      assign  SLAVE_RUSER[(6+1)*USER_WIDTH-1:6*USER_WIDTH]                                     = SLAVE6_RUSER;  
      assign  SLAVE_RVALID[6]                                                                  = SLAVE6_RVALID;
    end
      
  if ( NUM_SLAVES > 7 )
    begin
      //===================================================================
      //Slave7 Combine Signals
      //===================================================================
      //======================= SLAVE7 TO/FROM External Side=================
      //Outputs
      assign  SLAVE7_AWID     = SLAVE_AWID[(7+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:7*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE7_AWADDR   = SLAVE_AWADDR[(7+1)*ADDR_WIDTH-1:7*ADDR_WIDTH];  
      assign  SLAVE7_AWLEN    = SLAVE_AWLEN[(7+1)*8-1:7*8];  
      assign  SLAVE7_AWSIZE   = SLAVE_AWSIZE[(7+1)*3-1:7*3];  
      assign  SLAVE7_AWBURST  = SLAVE_AWBURST[(7+1)*2-1:7*2];  
      assign  SLAVE7_AWLOCK   = SLAVE_AWLOCK[(7+1)*2-1:7*2];  
      assign  SLAVE7_AWCACHE  = SLAVE_AWCACHE[(7+1)*4-1:7*4];  
      assign  SLAVE7_AWPROT   = SLAVE_AWPROT[(7+1)*3-1:7*3];  
      assign  SLAVE7_AWREGION = SLAVE_AWREGION[(7+1)*4-1:7*4];   
      assign  SLAVE7_AWQOS    = SLAVE_AWQOS[(7+1)*4-1:7*4];  
      assign  SLAVE7_AWUSER   = SLAVE_AWUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH];  
      assign  SLAVE7_AWVALID  = SLAVE_AWVALID[7];  
      assign  SLAVE7_WID      = SLAVE_WID[(7+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:7*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE7_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(7+1)*13-1:13*7]-1:SDW_LOWER_VEC[(7+1)*13-1:13*7]];  
      assign  SLAVE7_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(7+1)*13-1:13*7]/8-1:SDW_LOWER_VEC[(7+1)*13-1:13*7]/8];  
      assign  SLAVE7_WLAST    = SLAVE_WLAST[7];  
      assign  SLAVE7_WUSER    = SLAVE_WUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH];  
      assign  SLAVE7_WVALID   = SLAVE_WVALID[7];      
      assign  SLAVE7_BREADY   = SLAVE_BREADY[7];        
      assign  SLAVE7_ARID     = SLAVE_ARID[(7+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:7*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE7_ARADDR   = SLAVE_ARADDR[(7+1)*ADDR_WIDTH-1:7*ADDR_WIDTH];  
      assign  SLAVE7_ARLEN    = SLAVE_ARLEN[(7+1)*8-1:7*8];  
      assign  SLAVE7_ARSIZE   = SLAVE_ARSIZE[(7+1)*3-1:7*3];  
      assign  SLAVE7_ARBURST  = SLAVE_ARBURST[(7+1)*2-1:7*2];  
      assign  SLAVE7_ARLOCK   = SLAVE_ARLOCK[(7+1)*2-1:7*2];  
      assign  SLAVE7_ARCACHE  = SLAVE_ARCACHE[(7+1)*4-1:7*4] ;  
      assign  SLAVE7_ARPROT   = SLAVE_ARPROT[(7+1)*3-1:7*3] ;  
      assign  SLAVE7_ARREGION = SLAVE_ARREGION[(7+1)*4-1:7*4];   
      assign  SLAVE7_ARQOS    = SLAVE_ARQOS[(7+1)*4-1:7*4];  
      assign  SLAVE7_ARUSER   = SLAVE_ARUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH];  
      assign  SLAVE7_ARVALID  = SLAVE_ARVALID[7];      
      assign  SLAVE7_RREADY   = SLAVE_RREADY[7];  

      //Inputs      
      assign  SLAVE_AWREADY[7]                                                                 = SLAVE7_AWREADY;          
      assign  SLAVE_WREADY[7]                                                                  = SLAVE7_WREADY;        
      assign  SLAVE_BID[(7+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:7*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE7_BID;  
      assign  SLAVE_BRESP[(7+1)*2-1:7*2]                                                       = SLAVE7_BRESP;  
      assign  SLAVE_BUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH]                                     = SLAVE7_BUSER;  
      assign  SLAVE_BVALID[7]                                                                  = SLAVE7_BVALID;        
      assign  SLAVE_ARREADY[7]                                                                 = SLAVE7_ARREADY;        
      assign  SLAVE_RID[(7+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:7*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE7_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(7+1)*13-1:13*7]-1:SDW_LOWER_VEC[(7+1)*13-1:13*7]]     = SLAVE7_RDATA;  
      assign  SLAVE_RRESP[(7+1)*2-1:7*2]                                                       = SLAVE7_RRESP;  
      assign  SLAVE_RLAST[7]                                                                   = SLAVE7_RLAST;  
      assign  SLAVE_RUSER[(7+1)*USER_WIDTH-1:7*USER_WIDTH]                                     = SLAVE7_RUSER;  
      assign  SLAVE_RVALID[7]                                                                  = SLAVE7_RVALID;
    end
    
   
    
    if ( NUM_SLAVES > 8 )
    begin
      //===================================================================
      //Slave8 Combine Signals
      //===================================================================
      //======================= SLAVE8 TO/FROM External Side=================
      //Outputs
      assign  SLAVE8_AWID     = SLAVE_AWID[(8+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:8*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE8_AWADDR   = SLAVE_AWADDR[(8+1)*ADDR_WIDTH-1:8*ADDR_WIDTH];  
      assign  SLAVE8_AWLEN    = SLAVE_AWLEN[(8+1)*8-1:8*8];  
      assign  SLAVE8_AWSIZE   = SLAVE_AWSIZE[(8+1)*3-1:8*3];  
      assign  SLAVE8_AWBURST  = SLAVE_AWBURST[(8+1)*2-1:8*2];  
      assign  SLAVE8_AWLOCK   = SLAVE_AWLOCK[(8+1)*2-1:8*2];  
      assign  SLAVE8_AWCACHE  = SLAVE_AWCACHE[(8+1)*4-1:8*4];  
      assign  SLAVE8_AWPROT   = SLAVE_AWPROT[(8+1)*3-1:8*3];  
      assign  SLAVE8_AWREGION = SLAVE_AWREGION[(8+1)*4-1:8*4];   
      assign  SLAVE8_AWQOS    = SLAVE_AWQOS[(8+1)*4-1:8*4];  
      assign  SLAVE8_AWUSER   = SLAVE_AWUSER[(8+1)*USER_WIDTH-1:8*USER_WIDTH];  
      assign  SLAVE8_AWVALID  = SLAVE_AWVALID[8];  
      assign  SLAVE8_WID      = SLAVE_WID[(8+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:8*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE8_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(8+1)*13-1:13*8]-1:SDW_LOWER_VEC[(8+1)*13-1:13*8]];  
      assign  SLAVE8_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(8+1)*13-1:13*8]/8-1:SDW_LOWER_VEC[(8+1)*13-1:13*8]/8];  
      assign  SLAVE8_WLAST    = SLAVE_WLAST[8];  
      assign  SLAVE8_WUSER    = SLAVE_WUSER[(8+1)*USER_WIDTH-1:8*USER_WIDTH];  
      assign  SLAVE8_WVALID   = SLAVE_WVALID[8];      
      assign  SLAVE8_BREADY   = SLAVE_BREADY[8];        
      assign  SLAVE8_ARID     = SLAVE_ARID[(8+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:8*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE8_ARADDR   = SLAVE_ARADDR[(8+1)*ADDR_WIDTH-1:8*ADDR_WIDTH];  
      assign  SLAVE8_ARLEN    = SLAVE_ARLEN[(8+1)*8-1:8*8];  
      assign  SLAVE8_ARSIZE   = SLAVE_ARSIZE[(8+1)*3-1:8*3];  
      assign  SLAVE8_ARBURST  = SLAVE_ARBURST[(8+1)*2-1:8*2];  
      assign  SLAVE8_ARLOCK   = SLAVE_ARLOCK[(8+1)*2-1:8*2];  
      assign  SLAVE8_ARCACHE  = SLAVE_ARCACHE[(8+1)*4-1:8*4] ;  
      assign  SLAVE8_ARPROT   = SLAVE_ARPROT[(8+1)*3-1:8*3] ;  
      assign  SLAVE8_ARREGION = SLAVE_ARREGION[(8+1)*4-1:8*4];   
      assign  SLAVE8_ARQOS    = SLAVE_ARQOS[(8+1)*4-1:8*4];  
      assign  SLAVE8_ARUSER   = SLAVE_ARUSER[(8+1)*USER_WIDTH-1:8*USER_WIDTH];  
      assign  SLAVE8_ARVALID  = SLAVE_ARVALID[8];      
      assign  SLAVE8_RREADY   = SLAVE_RREADY[8];  

      //Inputs      
      assign  SLAVE_AWREADY[8]                                                                 = SLAVE8_AWREADY;          
      assign  SLAVE_WREADY[8]                                                                  = SLAVE8_WREADY;        
      assign  SLAVE_BID[(8+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:8*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE8_BID;  
      assign  SLAVE_BRESP[(8+1)*2-1:8*2]                                                       = SLAVE8_BRESP;  
      assign  SLAVE_BUSER[(8+1)*USER_WIDTH-1:8*USER_WIDTH]                                     = SLAVE8_BUSER;  
      assign  SLAVE_BVALID[8]                                                                  = SLAVE8_BVALID;        
      assign  SLAVE_ARREADY[8]                                                                 = SLAVE8_ARREADY;        
      assign  SLAVE_RID[(8+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:8*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE8_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(8+1)*13-1:13*8]-1:SDW_LOWER_VEC[(8+1)*13-1:13*8]]     = SLAVE8_RDATA;  
      assign  SLAVE_RRESP[(8+1)*2-1:8*2]                                                       = SLAVE8_RRESP;  
      assign  SLAVE_RLAST[8]                                                                   = SLAVE8_RLAST;  
      assign  SLAVE_RUSER[(8+1)*USER_WIDTH-1:8*USER_WIDTH]                                     = SLAVE8_RUSER;  
      assign  SLAVE_RVALID[8]                                                                  = SLAVE8_RVALID;
    end
    
    if ( NUM_SLAVES > 9 )
    begin
      //===================================================================
      //Slave9 Combine Signals
      //===================================================================
      //======================= SLAVE9 TO/FROM External Side=================
      //Outputs
      assign  SLAVE9_AWID     = SLAVE_AWID[(9+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:9*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE9_AWADDR   = SLAVE_AWADDR[(9+1)*ADDR_WIDTH-1:9*ADDR_WIDTH];  
      assign  SLAVE9_AWLEN    = SLAVE_AWLEN[(9+1)*8-1:9*8];  
      assign  SLAVE9_AWSIZE   = SLAVE_AWSIZE[(9+1)*3-1:9*3];  
      assign  SLAVE9_AWBURST  = SLAVE_AWBURST[(9+1)*2-1:9*2];  
      assign  SLAVE9_AWLOCK   = SLAVE_AWLOCK[(9+1)*2-1:9*2];  
      assign  SLAVE9_AWCACHE  = SLAVE_AWCACHE[(9+1)*4-1:9*4];  
      assign  SLAVE9_AWPROT   = SLAVE_AWPROT[(9+1)*3-1:9*3];  
      assign  SLAVE9_AWREGION = SLAVE_AWREGION[(9+1)*4-1:9*4];   
      assign  SLAVE9_AWQOS    = SLAVE_AWQOS[(9+1)*4-1:9*4];  
      assign  SLAVE9_AWUSER   = SLAVE_AWUSER[(9+1)*USER_WIDTH-1:9*USER_WIDTH];  
      assign  SLAVE9_AWVALID  = SLAVE_AWVALID[9];  
      assign  SLAVE9_WID      = SLAVE_WID[(9+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:9*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE9_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(9+1)*13-1:13*9]-1:SDW_LOWER_VEC[(9+1)*13-1:13*9]];  
      assign  SLAVE9_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(9+1)*13-1:13*9]/8-1:SDW_LOWER_VEC[(9+1)*13-1:13*9]/8];  
      assign  SLAVE9_WLAST    = SLAVE_WLAST[9];  
      assign  SLAVE9_WUSER    = SLAVE_WUSER[(9+1)*USER_WIDTH-1:9*USER_WIDTH];  
      assign  SLAVE9_WVALID   = SLAVE_WVALID[9];      
      assign  SLAVE9_BREADY   = SLAVE_BREADY[9];        
      assign  SLAVE9_ARID     = SLAVE_ARID[(9+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:9*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE9_ARADDR   = SLAVE_ARADDR[(9+1)*ADDR_WIDTH-1:9*ADDR_WIDTH];  
      assign  SLAVE9_ARLEN    = SLAVE_ARLEN[(9+1)*8-1:9*8];  
      assign  SLAVE9_ARSIZE   = SLAVE_ARSIZE[(9+1)*3-1:9*3];  
      assign  SLAVE9_ARBURST  = SLAVE_ARBURST[(9+1)*2-1:9*2];  
      assign  SLAVE9_ARLOCK   = SLAVE_ARLOCK[(9+1)*2-1:9*2];  
      assign  SLAVE9_ARCACHE  = SLAVE_ARCACHE[(9+1)*4-1:9*4] ;  
      assign  SLAVE9_ARPROT   = SLAVE_ARPROT[(9+1)*3-1:9*3] ;  
      assign  SLAVE9_ARREGION = SLAVE_ARREGION[(9+1)*4-1:9*4];   
      assign  SLAVE9_ARQOS    = SLAVE_ARQOS[(9+1)*4-1:9*4];  
      assign  SLAVE9_ARUSER   = SLAVE_ARUSER[(9+1)*USER_WIDTH-1:9*USER_WIDTH];  
      assign  SLAVE9_ARVALID  = SLAVE_ARVALID[9];      
      assign  SLAVE9_RREADY   = SLAVE_RREADY[9];  

      //Inputs      
      assign  SLAVE_AWREADY[9]                                                                 = SLAVE9_AWREADY;          
      assign  SLAVE_WREADY[9]                                                                  = SLAVE9_WREADY;        
      assign  SLAVE_BID[(9+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:9*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE9_BID;  
      assign  SLAVE_BRESP[(9+1)*2-1:9*2]                                                       = SLAVE9_BRESP;  
      assign  SLAVE_BUSER[(9+1)*USER_WIDTH-1:9*USER_WIDTH]                                     = SLAVE9_BUSER;  
      assign  SLAVE_BVALID[9]                                                                  = SLAVE9_BVALID;        
      assign  SLAVE_ARREADY[9]                                                                 = SLAVE9_ARREADY;        
      assign  SLAVE_RID[(9+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:9*(NUM_MASTERS_WIDTH+ID_WIDTH)]   = SLAVE9_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(9+1)*13-1:13*9]-1:SDW_LOWER_VEC[(9+1)*13-1:13*9]]     = SLAVE9_RDATA;  
      assign  SLAVE_RRESP[(9+1)*2-1:9*2]                                                       = SLAVE9_RRESP;  
      assign  SLAVE_RLAST[9]                                                                   = SLAVE9_RLAST;  
      assign  SLAVE_RUSER[(9+1)*USER_WIDTH-1:9*USER_WIDTH]                                     = SLAVE9_RUSER;  
      assign  SLAVE_RVALID[9]                                                                  = SLAVE9_RVALID;
    end
    
    if ( NUM_SLAVES > 10 )
    begin
      //===================================================================
      //Slave10 Combine Signals
      //===================================================================
      //======================= SLAVE10 TO/FROM External Side=================
      //Outputs
      assign  SLAVE10_AWID     = SLAVE_AWID[(10+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:10*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE10_AWADDR   = SLAVE_AWADDR[(10+1)*ADDR_WIDTH-1:10*ADDR_WIDTH];  
      assign  SLAVE10_AWLEN    = SLAVE_AWLEN[(10+1)*8-1:10*8];  
      assign  SLAVE10_AWSIZE   = SLAVE_AWSIZE[(10+1)*3-1:10*3];  
      assign  SLAVE10_AWBURST  = SLAVE_AWBURST[(10+1)*2-1:10*2];  
      assign  SLAVE10_AWLOCK   = SLAVE_AWLOCK[(10+1)*2-1:10*2];  
      assign  SLAVE10_AWCACHE  = SLAVE_AWCACHE[(10+1)*4-1:10*4];  
      assign  SLAVE10_AWPROT   = SLAVE_AWPROT[(10+1)*3-1:10*3];  
      assign  SLAVE10_AWREGION = SLAVE_AWREGION[(10+1)*4-1:10*4];   
      assign  SLAVE10_AWQOS    = SLAVE_AWQOS[(10+1)*4-1:10*4];  
      assign  SLAVE10_AWUSER   = SLAVE_AWUSER[(10+1)*USER_WIDTH-1:10*USER_WIDTH];  
      assign  SLAVE10_AWVALID  = SLAVE_AWVALID[10];  
      assign  SLAVE10_WID      = SLAVE_WID[(10+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:10*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE10_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(10+1)*13-1:13*10]-1:SDW_LOWER_VEC[(10+1)*13-1:13*10]];  
      assign  SLAVE10_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(10+1)*13-1:13*10]/8-1:SDW_LOWER_VEC[(10+1)*13-1:13*10]/8];  
      assign  SLAVE10_WLAST    = SLAVE_WLAST[10];  
      assign  SLAVE10_WUSER    = SLAVE_WUSER[(10+1)*USER_WIDTH-1:10*USER_WIDTH];  
      assign  SLAVE10_WVALID   = SLAVE_WVALID[10];      
      assign  SLAVE10_BREADY   = SLAVE_BREADY[10];        
      assign  SLAVE10_ARID     = SLAVE_ARID[(10+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:10*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE10_ARADDR   = SLAVE_ARADDR[(10+1)*ADDR_WIDTH-1:10*ADDR_WIDTH];  
      assign  SLAVE10_ARLEN    = SLAVE_ARLEN[(10+1)*8-1:10*8];  
      assign  SLAVE10_ARSIZE   = SLAVE_ARSIZE[(10+1)*3-1:10*3];  
      assign  SLAVE10_ARBURST  = SLAVE_ARBURST[(10+1)*2-1:10*2];  
      assign  SLAVE10_ARLOCK   = SLAVE_ARLOCK[(10+1)*2-1:10*2];  
      assign  SLAVE10_ARCACHE  = SLAVE_ARCACHE[(10+1)*4-1:10*4] ;  
      assign  SLAVE10_ARPROT   = SLAVE_ARPROT[(10+1)*3-1:10*3] ;  
      assign  SLAVE10_ARREGION = SLAVE_ARREGION[(10+1)*4-1:10*4];   
      assign  SLAVE10_ARQOS    = SLAVE_ARQOS[(10+1)*4-1:10*4];  
      assign  SLAVE10_ARUSER   = SLAVE_ARUSER[(10+1)*USER_WIDTH-1:10*USER_WIDTH];  
      assign  SLAVE10_ARVALID  = SLAVE_ARVALID[10];      
      assign  SLAVE10_RREADY   = SLAVE_RREADY[10];  

      //Inputs      
      assign  SLAVE_AWREADY[10]                                                                    = SLAVE10_AWREADY;          
      assign  SLAVE_WREADY[10]                                                                     = SLAVE10_WREADY;        
      assign  SLAVE_BID[(10+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:10*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE10_BID;  
      assign  SLAVE_BRESP[(10+1)*2-1:10*2]                                                         = SLAVE10_BRESP;  
      assign  SLAVE_BUSER[(10+1)*USER_WIDTH-1:10*USER_WIDTH]                                       = SLAVE10_BUSER;  
      assign  SLAVE_BVALID[10]                                                                     = SLAVE10_BVALID;        
      assign  SLAVE_ARREADY[10]                                                                    = SLAVE10_ARREADY;        
      assign  SLAVE_RID[(10+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:10*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE10_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(10+1)*13-1:13*10]-1:SDW_LOWER_VEC[(10+1)*13-1:13*10]]     = SLAVE10_RDATA;  
      assign  SLAVE_RRESP[(10+1)*2-1:10*2]                                                         = SLAVE10_RRESP;  
      assign  SLAVE_RLAST[10]                                                                      = SLAVE10_RLAST;  
      assign  SLAVE_RUSER[(10+1)*USER_WIDTH-1:10*USER_WIDTH]                                       = SLAVE10_RUSER;  
      assign  SLAVE_RVALID[10]                                                                     = SLAVE10_RVALID;
    end
    
    if ( NUM_SLAVES > 11 )
    begin
      //===================================================================
      //Slave11 Combine Signals
      //===================================================================
      //======================= SLAVE11 TO/FROM External Side=================
      //Outputs
      assign  SLAVE11_AWID     = SLAVE_AWID[(11+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:11*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE11_AWADDR   = SLAVE_AWADDR[(11+1)*ADDR_WIDTH-1:11*ADDR_WIDTH];  
      assign  SLAVE11_AWLEN    = SLAVE_AWLEN[(11+1)*8-1:11*8];  
      assign  SLAVE11_AWSIZE   = SLAVE_AWSIZE[(11+1)*3-1:11*3];  
      assign  SLAVE11_AWBURST  = SLAVE_AWBURST[(11+1)*2-1:11*2];  
      assign  SLAVE11_AWLOCK   = SLAVE_AWLOCK[(11+1)*2-1:11*2];  
      assign  SLAVE11_AWCACHE  = SLAVE_AWCACHE[(11+1)*4-1:11*4];  
      assign  SLAVE11_AWPROT   = SLAVE_AWPROT[(11+1)*3-1:11*3];  
      assign  SLAVE11_AWREGION = SLAVE_AWREGION[(11+1)*4-1:11*4];   
      assign  SLAVE11_AWQOS    = SLAVE_AWQOS[(11+1)*4-1:11*4];  
      assign  SLAVE11_AWUSER   = SLAVE_AWUSER[(11+1)*USER_WIDTH-1:11*USER_WIDTH];  
      assign  SLAVE11_AWVALID  = SLAVE_AWVALID[11];  
      assign  SLAVE11_WID      = SLAVE_WID[(11+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:11*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE11_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(11+1)*13-1:13*11]-1:SDW_LOWER_VEC[(11+1)*13-1:13*11]];  
      assign  SLAVE11_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(11+1)*13-1:13*11]/8-1:SDW_LOWER_VEC[(11+1)*13-1:13*11]/8];  
      assign  SLAVE11_WLAST    = SLAVE_WLAST[11];  
      assign  SLAVE11_WUSER    = SLAVE_WUSER[(11+1)*USER_WIDTH-1:11*USER_WIDTH];  
      assign  SLAVE11_WVALID   = SLAVE_WVALID[11];      
      assign  SLAVE11_BREADY   = SLAVE_BREADY[11];        
      assign  SLAVE11_ARID     = SLAVE_ARID[(11+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:11*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE11_ARADDR   = SLAVE_ARADDR[(11+1)*ADDR_WIDTH-1:11*ADDR_WIDTH];  
      assign  SLAVE11_ARLEN    = SLAVE_ARLEN[(11+1)*8-1:11*8];  
      assign  SLAVE11_ARSIZE   = SLAVE_ARSIZE[(11+1)*3-1:11*3];  
      assign  SLAVE11_ARBURST  = SLAVE_ARBURST[(11+1)*2-1:11*2];  
      assign  SLAVE11_ARLOCK   = SLAVE_ARLOCK[(11+1)*2-1:11*2];  
      assign  SLAVE11_ARCACHE  = SLAVE_ARCACHE[(11+1)*4-1:11*4] ;  
      assign  SLAVE11_ARPROT   = SLAVE_ARPROT[(11+1)*3-1:11*3] ;  
      assign  SLAVE11_ARREGION = SLAVE_ARREGION[(11+1)*4-1:11*4];   
      assign  SLAVE11_ARQOS    = SLAVE_ARQOS[(11+1)*4-1:11*4];  
      assign  SLAVE11_ARUSER   = SLAVE_ARUSER[(11+1)*USER_WIDTH-1:11*USER_WIDTH];  
      assign  SLAVE11_ARVALID  = SLAVE_ARVALID[11];      
      assign  SLAVE11_RREADY   = SLAVE_RREADY[11];  

      //Inputs      
      assign  SLAVE_AWREADY[11]                                                                    = SLAVE11_AWREADY;          
      assign  SLAVE_WREADY[11]                                                                     = SLAVE11_WREADY;        
      assign  SLAVE_BID[(11+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:11*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE11_BID;  
      assign  SLAVE_BRESP[(11+1)*2-1:11*2]                                                         = SLAVE11_BRESP;  
      assign  SLAVE_BUSER[(11+1)*USER_WIDTH-1:11*USER_WIDTH]                                       = SLAVE11_BUSER;  
      assign  SLAVE_BVALID[11]                                                                     = SLAVE11_BVALID;        
      assign  SLAVE_ARREADY[11]                                                                    = SLAVE11_ARREADY;        
      assign  SLAVE_RID[(11+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:11*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE11_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(11+1)*13-1:13*11]-1:SDW_LOWER_VEC[(11+1)*13-1:13*11]]     = SLAVE11_RDATA;  
      assign  SLAVE_RRESP[(11+1)*2-1:11*2]                                                         = SLAVE11_RRESP;  
      assign  SLAVE_RLAST[11]                                                                      = SLAVE11_RLAST;  
      assign  SLAVE_RUSER[(11+1)*USER_WIDTH-1:11*USER_WIDTH]                                       = SLAVE11_RUSER;  
      assign  SLAVE_RVALID[11]                                                                     = SLAVE11_RVALID;
    end
    
    if ( NUM_SLAVES > 12 )
    begin
      //===================================================================
      //Slave12 Combine Signals
      //===================================================================
      //======================= SLAVE12 TO/FROM External Side=================
      //Outputs
      assign  SLAVE12_AWID     = SLAVE_AWID[(12+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:12*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE12_AWADDR   = SLAVE_AWADDR[(12+1)*ADDR_WIDTH-1:12*ADDR_WIDTH];  
      assign  SLAVE12_AWLEN    = SLAVE_AWLEN[(12+1)*8-1:12*8];  
      assign  SLAVE12_AWSIZE   = SLAVE_AWSIZE[(12+1)*3-1:12*3];  
      assign  SLAVE12_AWBURST  = SLAVE_AWBURST[(12+1)*2-1:12*2];  
      assign  SLAVE12_AWLOCK   = SLAVE_AWLOCK[(12+1)*2-1:12*2];  
      assign  SLAVE12_AWCACHE  = SLAVE_AWCACHE[(12+1)*4-1:12*4];  
      assign  SLAVE12_AWPROT   = SLAVE_AWPROT[(12+1)*3-1:12*3];  
      assign  SLAVE12_AWREGION = SLAVE_AWREGION[(12+1)*4-1:12*4];   
      assign  SLAVE12_AWQOS    = SLAVE_AWQOS[(12+1)*4-1:12*4];  
      assign  SLAVE12_AWUSER   = SLAVE_AWUSER[(12+1)*USER_WIDTH-1:12*USER_WIDTH];  
      assign  SLAVE12_AWVALID  = SLAVE_AWVALID[12];  
      assign  SLAVE12_WID      = SLAVE_WID[(12+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:12*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE12_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(12+1)*13-1:13*12]-1:SDW_LOWER_VEC[(12+1)*13-1:13*12]];  
      assign  SLAVE12_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(12+1)*13-1:13*12]/8-1:SDW_LOWER_VEC[(12+1)*13-1:13*12]/8];  
      assign  SLAVE12_WLAST    = SLAVE_WLAST[12];  
      assign  SLAVE12_WUSER    = SLAVE_WUSER[(12+1)*USER_WIDTH-1:12*USER_WIDTH];  
      assign  SLAVE12_WVALID   = SLAVE_WVALID[12];      
      assign  SLAVE12_BREADY   = SLAVE_BREADY[12];        
      assign  SLAVE12_ARID     = SLAVE_ARID[(12+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:12*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE12_ARADDR   = SLAVE_ARADDR[(12+1)*ADDR_WIDTH-1:12*ADDR_WIDTH];  
      assign  SLAVE12_ARLEN    = SLAVE_ARLEN[(12+1)*8-1:12*8];  
      assign  SLAVE12_ARSIZE   = SLAVE_ARSIZE[(12+1)*3-1:12*3];  
      assign  SLAVE12_ARBURST  = SLAVE_ARBURST[(12+1)*2-1:12*2];  
      assign  SLAVE12_ARLOCK   = SLAVE_ARLOCK[(12+1)*2-1:12*2];  
      assign  SLAVE12_ARCACHE  = SLAVE_ARCACHE[(12+1)*4-1:12*4] ;  
      assign  SLAVE12_ARPROT   = SLAVE_ARPROT[(12+1)*3-1:12*3] ;  
      assign  SLAVE12_ARREGION = SLAVE_ARREGION[(12+1)*4-1:12*4];   
      assign  SLAVE12_ARQOS    = SLAVE_ARQOS[(12+1)*4-1:12*4];  
      assign  SLAVE12_ARUSER   = SLAVE_ARUSER[(12+1)*USER_WIDTH-1:12*USER_WIDTH];  
      assign  SLAVE12_ARVALID  = SLAVE_ARVALID[12];      
      assign  SLAVE12_RREADY   = SLAVE_RREADY[12];  

      //Inputs      
      assign  SLAVE_AWREADY[12]                                                                    = SLAVE12_AWREADY;          
      assign  SLAVE_WREADY[12]                                                                     = SLAVE12_WREADY;        
      assign  SLAVE_BID[(12+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:12*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE12_BID;  
      assign  SLAVE_BRESP[(12+1)*2-1:12*2]                                                         = SLAVE12_BRESP;  
      assign  SLAVE_BUSER[(12+1)*USER_WIDTH-1:12*USER_WIDTH]                                       = SLAVE12_BUSER;  
      assign  SLAVE_BVALID[12]                                                                     = SLAVE12_BVALID;        
      assign  SLAVE_ARREADY[12]                                                                    = SLAVE12_ARREADY;        
      assign  SLAVE_RID[(12+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:12*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE12_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(12+1)*13-1:13*12]-1:SDW_LOWER_VEC[(12+1)*13-1:13*12]]     = SLAVE12_RDATA;  
      assign  SLAVE_RRESP[(12+1)*2-1:12*2]                                                         = SLAVE12_RRESP;  
      assign  SLAVE_RLAST[12]                                                                      = SLAVE12_RLAST;  
      assign  SLAVE_RUSER[(12+1)*USER_WIDTH-1:12*USER_WIDTH]                                       = SLAVE12_RUSER;  
      assign  SLAVE_RVALID[12]                                                                     = SLAVE12_RVALID;
    end
    
    if ( NUM_SLAVES > 13 )
    begin
      //===================================================================
      //Slave13 Combine Signals
      //===================================================================
      //======================= SLAVE13 TO/FROM External Side=================
      //Outputs
      assign  SLAVE13_AWID     = SLAVE_AWID[(13+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:13*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE13_AWADDR   = SLAVE_AWADDR[(13+1)*ADDR_WIDTH-1:13*ADDR_WIDTH];  
      assign  SLAVE13_AWLEN    = SLAVE_AWLEN[(13+1)*8-1:13*8];  
      assign  SLAVE13_AWSIZE   = SLAVE_AWSIZE[(13+1)*3-1:13*3];  
      assign  SLAVE13_AWBURST  = SLAVE_AWBURST[(13+1)*2-1:13*2];  
      assign  SLAVE13_AWLOCK   = SLAVE_AWLOCK[(13+1)*2-1:13*2];  
      assign  SLAVE13_AWCACHE  = SLAVE_AWCACHE[(13+1)*4-1:13*4];  
      assign  SLAVE13_AWPROT   = SLAVE_AWPROT[(13+1)*3-1:13*3];  
      assign  SLAVE13_AWREGION = SLAVE_AWREGION[(13+1)*4-1:13*4];   
      assign  SLAVE13_AWQOS    = SLAVE_AWQOS[(13+1)*4-1:13*4];  
      assign  SLAVE13_AWUSER   = SLAVE_AWUSER[(13+1)*USER_WIDTH-1:13*USER_WIDTH];  
      assign  SLAVE13_AWVALID  = SLAVE_AWVALID[13];  
      assign  SLAVE13_WID      = SLAVE_WID[(13+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:13*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE13_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(13+1)*13-1:13*13]-1:SDW_LOWER_VEC[(13+1)*13-1:13*13]];  
      assign  SLAVE13_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(13+1)*13-1:13*13]/8-1:SDW_LOWER_VEC[(13+1)*13-1:13*13]/8];  
      assign  SLAVE13_WLAST    = SLAVE_WLAST[13];  
      assign  SLAVE13_WUSER    = SLAVE_WUSER[(13+1)*USER_WIDTH-1:13*USER_WIDTH];  
      assign  SLAVE13_WVALID   = SLAVE_WVALID[13];      
      assign  SLAVE13_BREADY   = SLAVE_BREADY[13];        
      assign  SLAVE13_ARID     = SLAVE_ARID[(13+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:13*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE13_ARADDR   = SLAVE_ARADDR[(13+1)*ADDR_WIDTH-1:13*ADDR_WIDTH];  
      assign  SLAVE13_ARLEN    = SLAVE_ARLEN[(13+1)*8-1:13*8];  
      assign  SLAVE13_ARSIZE   = SLAVE_ARSIZE[(13+1)*3-1:13*3];  
      assign  SLAVE13_ARBURST  = SLAVE_ARBURST[(13+1)*2-1:13*2];  
      assign  SLAVE13_ARLOCK   = SLAVE_ARLOCK[(13+1)*2-1:13*2];  
      assign  SLAVE13_ARCACHE  = SLAVE_ARCACHE[(13+1)*4-1:13*4] ;  
      assign  SLAVE13_ARPROT   = SLAVE_ARPROT[(13+1)*3-1:13*3] ;  
      assign  SLAVE13_ARREGION = SLAVE_ARREGION[(13+1)*4-1:13*4];   
      assign  SLAVE13_ARQOS    = SLAVE_ARQOS[(13+1)*4-1:13*4];  
      assign  SLAVE13_ARUSER   = SLAVE_ARUSER[(13+1)*USER_WIDTH-1:13*USER_WIDTH];  
      assign  SLAVE13_ARVALID  = SLAVE_ARVALID[13];      
      assign  SLAVE13_RREADY   = SLAVE_RREADY[13];  

      //Inputs      
      assign  SLAVE_AWREADY[13]                                                                    = SLAVE13_AWREADY;          
      assign  SLAVE_WREADY[13]                                                                     = SLAVE13_WREADY;        
      assign  SLAVE_BID[(13+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:13*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE13_BID;  
      assign  SLAVE_BRESP[(13+1)*2-1:13*2]                                                         = SLAVE13_BRESP;  
      assign  SLAVE_BUSER[(13+1)*USER_WIDTH-1:13*USER_WIDTH]                                       = SLAVE13_BUSER;  
      assign  SLAVE_BVALID[13]                                                                     = SLAVE13_BVALID;        
      assign  SLAVE_ARREADY[13]                                                                    = SLAVE13_ARREADY;        
      assign  SLAVE_RID[(13+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:13*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE13_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(13+1)*13-1:13*13]-1:SDW_LOWER_VEC[(13+1)*13-1:13*13]]     = SLAVE13_RDATA;  
      assign  SLAVE_RRESP[(13+1)*2-1:13*2]                                                         = SLAVE13_RRESP;  
      assign  SLAVE_RLAST[13]                                                                      = SLAVE13_RLAST;  
      assign  SLAVE_RUSER[(13+1)*USER_WIDTH-1:13*USER_WIDTH]                                       = SLAVE13_RUSER;  
      assign  SLAVE_RVALID[13]                                                                     = SLAVE13_RVALID;
    end
    
    if ( NUM_SLAVES > 14 )
    begin
      //===================================================================
      //Slave14 Combine Signals
      //===================================================================
      //======================= SLAVE14 TO/FROM External Side=================
      //Outputs
      assign  SLAVE14_AWID     = SLAVE_AWID[(14+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:14*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE14_AWADDR   = SLAVE_AWADDR[(14+1)*ADDR_WIDTH-1:14*ADDR_WIDTH];  
      assign  SLAVE14_AWLEN    = SLAVE_AWLEN[(14+1)*8-1:14*8];  
      assign  SLAVE14_AWSIZE   = SLAVE_AWSIZE[(14+1)*3-1:14*3];  
      assign  SLAVE14_AWBURST  = SLAVE_AWBURST[(14+1)*2-1:14*2];  
      assign  SLAVE14_AWLOCK   = SLAVE_AWLOCK[(14+1)*2-1:14*2];  
      assign  SLAVE14_AWCACHE  = SLAVE_AWCACHE[(14+1)*4-1:14*4];  
      assign  SLAVE14_AWPROT   = SLAVE_AWPROT[(14+1)*3-1:14*3];  
      assign  SLAVE14_AWREGION = SLAVE_AWREGION[(14+1)*4-1:14*4];   
      assign  SLAVE14_AWQOS    = SLAVE_AWQOS[(14+1)*4-1:14*4];  
      assign  SLAVE14_AWUSER   = SLAVE_AWUSER[(14+1)*USER_WIDTH-1:14*USER_WIDTH];  
      assign  SLAVE14_AWVALID  = SLAVE_AWVALID[14];  
      assign  SLAVE14_WID      = SLAVE_WID[(14+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:14*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE14_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(14+1)*13-1:13*14]-1:SDW_LOWER_VEC[(14+1)*13-1:13*14]];  
      assign  SLAVE14_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(14+1)*13-1:13*14]/8-1:SDW_LOWER_VEC[(14+1)*13-1:13*14]/8];  
      assign  SLAVE14_WLAST    = SLAVE_WLAST[14];  
      assign  SLAVE14_WUSER    = SLAVE_WUSER[(14+1)*USER_WIDTH-1:14*USER_WIDTH];  
      assign  SLAVE14_WVALID   = SLAVE_WVALID[14];      
      assign  SLAVE14_BREADY   = SLAVE_BREADY[14];        
      assign  SLAVE14_ARID     = SLAVE_ARID[(14+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:14*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE14_ARADDR   = SLAVE_ARADDR[(14+1)*ADDR_WIDTH-1:14*ADDR_WIDTH];  
      assign  SLAVE14_ARLEN    = SLAVE_ARLEN[(14+1)*8-1:14*8];  
      assign  SLAVE14_ARSIZE   = SLAVE_ARSIZE[(14+1)*3-1:14*3];  
      assign  SLAVE14_ARBURST  = SLAVE_ARBURST[(14+1)*2-1:14*2];  
      assign  SLAVE14_ARLOCK   = SLAVE_ARLOCK[(14+1)*2-1:14*2];  
      assign  SLAVE14_ARCACHE  = SLAVE_ARCACHE[(14+1)*4-1:14*4] ;  
      assign  SLAVE14_ARPROT   = SLAVE_ARPROT[(14+1)*3-1:14*3] ;  
      assign  SLAVE14_ARREGION = SLAVE_ARREGION[(14+1)*4-1:14*4];   
      assign  SLAVE14_ARQOS    = SLAVE_ARQOS[(14+1)*4-1:14*4];  
      assign  SLAVE14_ARUSER   = SLAVE_ARUSER[(14+1)*USER_WIDTH-1:14*USER_WIDTH];  
      assign  SLAVE14_ARVALID  = SLAVE_ARVALID[14];      
      assign  SLAVE14_RREADY   = SLAVE_RREADY[14];  

      //Inputs      
      assign  SLAVE_AWREADY[14]                                                                    = SLAVE14_AWREADY;
      assign  SLAVE_WREADY[14]                                                                     = SLAVE14_WREADY;
      assign  SLAVE_BID[(14+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:14*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE14_BID;
      assign  SLAVE_BRESP[(14+1)*2-1:14*2]                                                         = SLAVE14_BRESP;
      assign  SLAVE_BUSER[(14+1)*USER_WIDTH-1:14*USER_WIDTH]                                       = SLAVE14_BUSER;
      assign  SLAVE_BVALID[14]                                                                     = SLAVE14_BVALID;
      assign  SLAVE_ARREADY[14]                                                                    = SLAVE14_ARREADY;
      assign  SLAVE_RID[(14+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:14*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE14_RID;
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(14+1)*13-1:13*14]-1:SDW_LOWER_VEC[(14+1)*13-1:13*14]]     = SLAVE14_RDATA;
      assign  SLAVE_RRESP[(14+1)*2-1:14*2]                                                         = SLAVE14_RRESP;
      assign  SLAVE_RLAST[14]                                                                      = SLAVE14_RLAST;
      assign  SLAVE_RUSER[(14+1)*USER_WIDTH-1:14*USER_WIDTH]                                       = SLAVE14_RUSER;
      assign  SLAVE_RVALID[14]                                                                     = SLAVE14_RVALID;
    end
    
    if ( NUM_SLAVES > 15 )
    begin
      //===================================================================
      //Slave15 Combine Signals
      //===================================================================
      //======================= SLAVE15 TO/FROM External Side=================
      //Outputs
      assign  SLAVE15_AWID     = SLAVE_AWID[(15+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:15*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE15_AWADDR   = SLAVE_AWADDR[(15+1)*ADDR_WIDTH-1:15*ADDR_WIDTH];  
      assign  SLAVE15_AWLEN    = SLAVE_AWLEN[(15+1)*8-1:15*8];  
      assign  SLAVE15_AWSIZE   = SLAVE_AWSIZE[(15+1)*3-1:15*3];  
      assign  SLAVE15_AWBURST  = SLAVE_AWBURST[(15+1)*2-1:15*2];  
      assign  SLAVE15_AWLOCK   = SLAVE_AWLOCK[(15+1)*2-1:15*2];  
      assign  SLAVE15_AWCACHE  = SLAVE_AWCACHE[(15+1)*4-1:15*4];  
      assign  SLAVE15_AWPROT   = SLAVE_AWPROT[(15+1)*3-1:15*3];  
      assign  SLAVE15_AWREGION = SLAVE_AWREGION[(15+1)*4-1:15*4];   
      assign  SLAVE15_AWQOS    = SLAVE_AWQOS[(15+1)*4-1:15*4];  
      assign  SLAVE15_AWUSER   = SLAVE_AWUSER[(15+1)*USER_WIDTH-1:15*USER_WIDTH];  
      assign  SLAVE15_AWVALID  = SLAVE_AWVALID[15];  
      assign  SLAVE15_WID      = SLAVE_WID[(15+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:15*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE15_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(15+1)*13-1:13*15]-1:SDW_LOWER_VEC[(15+1)*13-1:13*15]];  
      assign  SLAVE15_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(15+1)*13-1:13*15]/8-1:SDW_LOWER_VEC[(15+1)*13-1:13*15]/8];  
      assign  SLAVE15_WLAST    = SLAVE_WLAST[15];  
      assign  SLAVE15_WUSER    = SLAVE_WUSER[(15+1)*USER_WIDTH-1:15*USER_WIDTH];  
      assign  SLAVE15_WVALID   = SLAVE_WVALID[15];      
      assign  SLAVE15_BREADY   = SLAVE_BREADY[15];        
      assign  SLAVE15_ARID     = SLAVE_ARID[(15+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:15*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE15_ARADDR   = SLAVE_ARADDR[(15+1)*ADDR_WIDTH-1:15*ADDR_WIDTH];  
      assign  SLAVE15_ARLEN    = SLAVE_ARLEN[(15+1)*8-1:15*8];  
      assign  SLAVE15_ARSIZE   = SLAVE_ARSIZE[(15+1)*3-1:15*3];  
      assign  SLAVE15_ARBURST  = SLAVE_ARBURST[(15+1)*2-1:15*2];  
      assign  SLAVE15_ARLOCK   = SLAVE_ARLOCK[(15+1)*2-1:15*2];  
      assign  SLAVE15_ARCACHE  = SLAVE_ARCACHE[(15+1)*4-1:15*4] ;  
      assign  SLAVE15_ARPROT   = SLAVE_ARPROT[(15+1)*3-1:15*3] ;  
      assign  SLAVE15_ARREGION = SLAVE_ARREGION[(15+1)*4-1:15*4];   
      assign  SLAVE15_ARQOS    = SLAVE_ARQOS[(15+1)*4-1:15*4];  
      assign  SLAVE15_ARUSER   = SLAVE_ARUSER[(15+1)*USER_WIDTH-1:15*USER_WIDTH];  
      assign  SLAVE15_ARVALID  = SLAVE_ARVALID[15];      
      assign  SLAVE15_RREADY   = SLAVE_RREADY[15];  

      //Inputs      
      assign  SLAVE_AWREADY[15]                                                                    = SLAVE15_AWREADY;          
      assign  SLAVE_WREADY[15]                                                                     = SLAVE15_WREADY;        
      assign  SLAVE_BID[(15+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:15*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE15_BID;  
      assign  SLAVE_BRESP[(15+1)*2-1:15*2]                                                         = SLAVE15_BRESP;  
      assign  SLAVE_BUSER[(15+1)*USER_WIDTH-1:15*USER_WIDTH]                                       = SLAVE15_BUSER;  
      assign  SLAVE_BVALID[15]                                                                     = SLAVE15_BVALID;        
      assign  SLAVE_ARREADY[15]                                                                    = SLAVE15_ARREADY;        
      assign  SLAVE_RID[(15+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:15*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE15_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(15+1)*13-1:13*15]-1:SDW_LOWER_VEC[(15+1)*13-1:13*15]]     = SLAVE15_RDATA;  
      assign  SLAVE_RRESP[(15+1)*2-1:15*2]                                                         = SLAVE15_RRESP;  
      assign  SLAVE_RLAST[15]                                                                      = SLAVE15_RLAST;  
      assign  SLAVE_RUSER[(15+1)*USER_WIDTH-1:15*USER_WIDTH]                                       = SLAVE15_RUSER;  
      assign  SLAVE_RVALID[15]                                                                     = SLAVE15_RVALID;
    end
    
    if ( NUM_SLAVES > 16 )
    begin
      //===================================================================
      //Slave16 Combine Signals
      //===================================================================
      //======================= SLAVE16 TO/FROM External Side=================
      //Outputs
      assign  SLAVE16_AWID     = SLAVE_AWID[(16+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:16*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE16_AWADDR   = SLAVE_AWADDR[(16+1)*ADDR_WIDTH-1:16*ADDR_WIDTH];  
      assign  SLAVE16_AWLEN    = SLAVE_AWLEN[(16+1)*8-1:16*8];  
      assign  SLAVE16_AWSIZE   = SLAVE_AWSIZE[(16+1)*3-1:16*3];  
      assign  SLAVE16_AWBURST  = SLAVE_AWBURST[(16+1)*2-1:16*2];  
      assign  SLAVE16_AWLOCK   = SLAVE_AWLOCK[(16+1)*2-1:16*2];  
      assign  SLAVE16_AWCACHE  = SLAVE_AWCACHE[(16+1)*4-1:16*4];  
      assign  SLAVE16_AWPROT   = SLAVE_AWPROT[(16+1)*3-1:16*3];  
      assign  SLAVE16_AWREGION = SLAVE_AWREGION[(16+1)*4-1:16*4];   
      assign  SLAVE16_AWQOS    = SLAVE_AWQOS[(16+1)*4-1:16*4];  
      assign  SLAVE16_AWUSER   = SLAVE_AWUSER[(16+1)*USER_WIDTH-1:16*USER_WIDTH];  
      assign  SLAVE16_AWVALID  = SLAVE_AWVALID[16];  
      assign  SLAVE16_WID      = SLAVE_WID[(16+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:16*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE16_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(16+1)*13-1:13*16]-1:SDW_LOWER_VEC[(16+1)*13-1:13*16]];  
      assign  SLAVE16_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(16+1)*13-1:13*16]/8-1:SDW_LOWER_VEC[(16+1)*13-1:13*16]/8];  
      assign  SLAVE16_WLAST    = SLAVE_WLAST[16];  
      assign  SLAVE16_WUSER    = SLAVE_WUSER[(16+1)*USER_WIDTH-1:16*USER_WIDTH];  
      assign  SLAVE16_WVALID   = SLAVE_WVALID[16];      
      assign  SLAVE16_BREADY   = SLAVE_BREADY[16];        
      assign  SLAVE16_ARID     = SLAVE_ARID[(16+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:16*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE16_ARADDR   = SLAVE_ARADDR[(16+1)*ADDR_WIDTH-1:16*ADDR_WIDTH];  
      assign  SLAVE16_ARLEN    = SLAVE_ARLEN[(16+1)*8-1:16*8];  
      assign  SLAVE16_ARSIZE   = SLAVE_ARSIZE[(16+1)*3-1:16*3];  
      assign  SLAVE16_ARBURST  = SLAVE_ARBURST[(16+1)*2-1:16*2];  
      assign  SLAVE16_ARLOCK   = SLAVE_ARLOCK[(16+1)*2-1:16*2];  
      assign  SLAVE16_ARCACHE  = SLAVE_ARCACHE[(16+1)*4-1:16*4] ;  
      assign  SLAVE16_ARPROT   = SLAVE_ARPROT[(16+1)*3-1:16*3] ;  
      assign  SLAVE16_ARREGION = SLAVE_ARREGION[(16+1)*4-1:16*4];   
      assign  SLAVE16_ARQOS    = SLAVE_ARQOS[(16+1)*4-1:16*4];  
      assign  SLAVE16_ARUSER   = SLAVE_ARUSER[(16+1)*USER_WIDTH-1:16*USER_WIDTH];  
      assign  SLAVE16_ARVALID  = SLAVE_ARVALID[16];      
      assign  SLAVE16_RREADY   = SLAVE_RREADY[16];  

      //Inputs      
      assign  SLAVE_AWREADY[16]                                                                    = SLAVE16_AWREADY;          
      assign  SLAVE_WREADY[16]                                                                     = SLAVE16_WREADY;        
      assign  SLAVE_BID[(16+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:16*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE16_BID;  
      assign  SLAVE_BRESP[(16+1)*2-1:16*2]                                                         = SLAVE16_BRESP;  
      assign  SLAVE_BUSER[(16+1)*USER_WIDTH-1:16*USER_WIDTH]                                       = SLAVE16_BUSER;  
      assign  SLAVE_BVALID[16]                                                                     = SLAVE16_BVALID;        
      assign  SLAVE_ARREADY[16]                                                                    = SLAVE16_ARREADY;        
      assign  SLAVE_RID[(16+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:16*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE16_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(16+1)*13-1:13*16]-1:SDW_LOWER_VEC[(16+1)*13-1:13*16]]     = SLAVE16_RDATA;  
      assign  SLAVE_RRESP[(16+1)*2-1:16*2]                                                         = SLAVE16_RRESP;  
      assign  SLAVE_RLAST[16]                                                                      = SLAVE16_RLAST;  
      assign  SLAVE_RUSER[(16+1)*USER_WIDTH-1:16*USER_WIDTH]                                       = SLAVE16_RUSER;  
      assign  SLAVE_RVALID[16]                                                                     = SLAVE16_RVALID;
    end
    
    if ( NUM_SLAVES > 17 )
    begin
      //===================================================================
      //Slave17 Combine Signals
      //===================================================================
      //======================= SLAVE17 TO/FROM External Side=================
      //Outputs
      assign  SLAVE17_AWID     = SLAVE_AWID[(17+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:17*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE17_AWADDR   = SLAVE_AWADDR[(17+1)*ADDR_WIDTH-1:17*ADDR_WIDTH];  
      assign  SLAVE17_AWLEN    = SLAVE_AWLEN[(17+1)*8-1:17*8];  
      assign  SLAVE17_AWSIZE   = SLAVE_AWSIZE[(17+1)*3-1:17*3];  
      assign  SLAVE17_AWBURST  = SLAVE_AWBURST[(17+1)*2-1:17*2];  
      assign  SLAVE17_AWLOCK   = SLAVE_AWLOCK[(17+1)*2-1:17*2];  
      assign  SLAVE17_AWCACHE  = SLAVE_AWCACHE[(17+1)*4-1:17*4];  
      assign  SLAVE17_AWPROT   = SLAVE_AWPROT[(17+1)*3-1:17*3];  
      assign  SLAVE17_AWREGION = SLAVE_AWREGION[(17+1)*4-1:17*4];   
      assign  SLAVE17_AWQOS    = SLAVE_AWQOS[(17+1)*4-1:17*4];  
      assign  SLAVE17_AWUSER   = SLAVE_AWUSER[(17+1)*USER_WIDTH-1:17*USER_WIDTH];  
      assign  SLAVE17_AWVALID  = SLAVE_AWVALID[17];  
      assign  SLAVE17_WID      = SLAVE_WID[(17+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:17*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE17_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(17+1)*13-1:13*17]-1:SDW_LOWER_VEC[(17+1)*13-1:13*17]];  
      assign  SLAVE17_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(17+1)*13-1:13*17]/8-1:SDW_LOWER_VEC[(17+1)*13-1:13*17]/8];  
      assign  SLAVE17_WLAST    = SLAVE_WLAST[17];  
      assign  SLAVE17_WUSER    = SLAVE_WUSER[(17+1)*USER_WIDTH-1:17*USER_WIDTH];  
      assign  SLAVE17_WVALID   = SLAVE_WVALID[17];      
      assign  SLAVE17_BREADY   = SLAVE_BREADY[17];        
      assign  SLAVE17_ARID     = SLAVE_ARID[(17+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:17*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE17_ARADDR   = SLAVE_ARADDR[(17+1)*ADDR_WIDTH-1:17*ADDR_WIDTH];  
      assign  SLAVE17_ARLEN    = SLAVE_ARLEN[(17+1)*8-1:17*8];  
      assign  SLAVE17_ARSIZE   = SLAVE_ARSIZE[(17+1)*3-1:17*3];  
      assign  SLAVE17_ARBURST  = SLAVE_ARBURST[(17+1)*2-1:17*2];  
      assign  SLAVE17_ARLOCK   = SLAVE_ARLOCK[(17+1)*2-1:17*2];  
      assign  SLAVE17_ARCACHE  = SLAVE_ARCACHE[(17+1)*4-1:17*4] ;  
      assign  SLAVE17_ARPROT   = SLAVE_ARPROT[(17+1)*3-1:17*3] ;  
      assign  SLAVE17_ARREGION = SLAVE_ARREGION[(17+1)*4-1:17*4];   
      assign  SLAVE17_ARQOS    = SLAVE_ARQOS[(17+1)*4-1:17*4];  
      assign  SLAVE17_ARUSER   = SLAVE_ARUSER[(17+1)*USER_WIDTH-1:17*USER_WIDTH];  
      assign  SLAVE17_ARVALID  = SLAVE_ARVALID[17];      
      assign  SLAVE17_RREADY   = SLAVE_RREADY[17];  

      //Inputs      
      assign  SLAVE_AWREADY[17]                                                                    = SLAVE17_AWREADY;          
      assign  SLAVE_WREADY[17]                                                                     = SLAVE17_WREADY;        
      assign  SLAVE_BID[(17+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:17*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE17_BID;  
      assign  SLAVE_BRESP[(17+1)*2-1:17*2]                                                         = SLAVE17_BRESP;  
      assign  SLAVE_BUSER[(17+1)*USER_WIDTH-1:17*USER_WIDTH]                                       = SLAVE17_BUSER;  
      assign  SLAVE_BVALID[17]                                                                     = SLAVE17_BVALID;        
      assign  SLAVE_ARREADY[17]                                                                    = SLAVE17_ARREADY;        
      assign  SLAVE_RID[(17+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:17*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE17_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(17+1)*13-1:13*17]-1:SDW_LOWER_VEC[(17+1)*13-1:13*17]]     = SLAVE17_RDATA;  
      assign  SLAVE_RRESP[(17+1)*2-1:17*2]                                                         = SLAVE17_RRESP;  
      assign  SLAVE_RLAST[17]                                                                      = SLAVE17_RLAST;  
      assign  SLAVE_RUSER[(17+1)*USER_WIDTH-1:17*USER_WIDTH]                                       = SLAVE17_RUSER;  
      assign  SLAVE_RVALID[17]                                                                     = SLAVE17_RVALID;
    end
    
    if ( NUM_SLAVES > 18 )
    begin
      //===================================================================
      //Slave18 Combine Signals
      //===================================================================
      //======================= SLAVE18 TO/FROM External Side=================
      //Outputs
      assign  SLAVE18_AWID     = SLAVE_AWID[(18+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:18*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE18_AWADDR   = SLAVE_AWADDR[(18+1)*ADDR_WIDTH-1:18*ADDR_WIDTH];  
      assign  SLAVE18_AWLEN    = SLAVE_AWLEN[(18+1)*8-1:18*8];  
      assign  SLAVE18_AWSIZE   = SLAVE_AWSIZE[(18+1)*3-1:18*3];  
      assign  SLAVE18_AWBURST  = SLAVE_AWBURST[(18+1)*2-1:18*2];  
      assign  SLAVE18_AWLOCK   = SLAVE_AWLOCK[(18+1)*2-1:18*2];  
      assign  SLAVE18_AWCACHE  = SLAVE_AWCACHE[(18+1)*4-1:18*4];  
      assign  SLAVE18_AWPROT   = SLAVE_AWPROT[(18+1)*3-1:18*3];  
      assign  SLAVE18_AWREGION = SLAVE_AWREGION[(18+1)*4-1:18*4];   
      assign  SLAVE18_AWQOS    = SLAVE_AWQOS[(18+1)*4-1:18*4];  
      assign  SLAVE18_AWUSER   = SLAVE_AWUSER[(18+1)*USER_WIDTH-1:18*USER_WIDTH];  
      assign  SLAVE18_AWVALID  = SLAVE_AWVALID[18];  
      assign  SLAVE18_WID      = SLAVE_WID[(18+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:18*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE18_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(18+1)*13-1:13*18]-1:SDW_LOWER_VEC[(18+1)*13-1:13*18]];  
      assign  SLAVE18_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(18+1)*13-1:13*18]/8-1:SDW_LOWER_VEC[(18+1)*13-1:13*18]/8];  
      assign  SLAVE18_WLAST    = SLAVE_WLAST[18];  
      assign  SLAVE18_WUSER    = SLAVE_WUSER[(18+1)*USER_WIDTH-1:18*USER_WIDTH];  
      assign  SLAVE18_WVALID   = SLAVE_WVALID[18];      
      assign  SLAVE18_BREADY   = SLAVE_BREADY[18];        
      assign  SLAVE18_ARID     = SLAVE_ARID[(18+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:18*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE18_ARADDR   = SLAVE_ARADDR[(18+1)*ADDR_WIDTH-1:18*ADDR_WIDTH];  
      assign  SLAVE18_ARLEN    = SLAVE_ARLEN[(18+1)*8-1:18*8];  
      assign  SLAVE18_ARSIZE   = SLAVE_ARSIZE[(18+1)*3-1:18*3];  
      assign  SLAVE18_ARBURST  = SLAVE_ARBURST[(18+1)*2-1:18*2];  
      assign  SLAVE18_ARLOCK   = SLAVE_ARLOCK[(18+1)*2-1:18*2];  
      assign  SLAVE18_ARCACHE  = SLAVE_ARCACHE[(18+1)*4-1:18*4] ;  
      assign  SLAVE18_ARPROT   = SLAVE_ARPROT[(18+1)*3-1:18*3] ;  
      assign  SLAVE18_ARREGION = SLAVE_ARREGION[(18+1)*4-1:18*4];   
      assign  SLAVE18_ARQOS    = SLAVE_ARQOS[(18+1)*4-1:18*4];  
      assign  SLAVE18_ARUSER   = SLAVE_ARUSER[(18+1)*USER_WIDTH-1:18*USER_WIDTH];  
      assign  SLAVE18_ARVALID  = SLAVE_ARVALID[18];      
      assign  SLAVE18_RREADY   = SLAVE_RREADY[18];  

      //Inputs      
      assign  SLAVE_AWREADY[18]                                                                    = SLAVE18_AWREADY;          
      assign  SLAVE_WREADY[18]                                                                     = SLAVE18_WREADY;        
      assign  SLAVE_BID[(18+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:18*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE18_BID;  
      assign  SLAVE_BRESP[(18+1)*2-1:18*2]                                                         = SLAVE18_BRESP;  
      assign  SLAVE_BUSER[(18+1)*USER_WIDTH-1:18*USER_WIDTH]                                       = SLAVE18_BUSER;  
      assign  SLAVE_BVALID[18]                                                                     = SLAVE18_BVALID;        
      assign  SLAVE_ARREADY[18]                                                                    = SLAVE18_ARREADY;        
      assign  SLAVE_RID[(18+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:18*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE18_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(18+1)*13-1:13*18]-1:SDW_LOWER_VEC[(18+1)*13-1:13*18]]     = SLAVE18_RDATA;  
      assign  SLAVE_RRESP[(18+1)*2-1:18*2]                                                         = SLAVE18_RRESP;  
      assign  SLAVE_RLAST[18]                                                                      = SLAVE18_RLAST;  
      assign  SLAVE_RUSER[(18+1)*USER_WIDTH-1:18*USER_WIDTH]                                       = SLAVE18_RUSER;  
      assign  SLAVE_RVALID[18]                                                                     = SLAVE18_RVALID;
    end
    
    if ( NUM_SLAVES > 19 )
    begin
      //===================================================================
      //Slave19 Combine Signals
      //===================================================================
      //======================= SLAVE19 TO/FROM External Side=================
      //Outputs
      assign  SLAVE19_AWID     = SLAVE_AWID[(19+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:19*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE19_AWADDR   = SLAVE_AWADDR[(19+1)*ADDR_WIDTH-1:19*ADDR_WIDTH];  
      assign  SLAVE19_AWLEN    = SLAVE_AWLEN[(19+1)*8-1:19*8];  
      assign  SLAVE19_AWSIZE   = SLAVE_AWSIZE[(19+1)*3-1:19*3];  
      assign  SLAVE19_AWBURST  = SLAVE_AWBURST[(19+1)*2-1:19*2];  
      assign  SLAVE19_AWLOCK   = SLAVE_AWLOCK[(19+1)*2-1:19*2];  
      assign  SLAVE19_AWCACHE  = SLAVE_AWCACHE[(19+1)*4-1:19*4];  
      assign  SLAVE19_AWPROT   = SLAVE_AWPROT[(19+1)*3-1:19*3];  
      assign  SLAVE19_AWREGION = SLAVE_AWREGION[(19+1)*4-1:19*4];   
      assign  SLAVE19_AWQOS    = SLAVE_AWQOS[(19+1)*4-1:19*4];  
      assign  SLAVE19_AWUSER   = SLAVE_AWUSER[(19+1)*USER_WIDTH-1:19*USER_WIDTH];  
      assign  SLAVE19_AWVALID  = SLAVE_AWVALID[19];  
      assign  SLAVE19_WID      = SLAVE_WID[(19+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:19*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE19_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(19+1)*13-1:13*19]-1:SDW_LOWER_VEC[(19+1)*13-1:13*19]];  
      assign  SLAVE19_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(19+1)*13-1:13*19]/8-1:SDW_LOWER_VEC[(19+1)*13-1:13*19]/8];  
      assign  SLAVE19_WLAST    = SLAVE_WLAST[19];  
      assign  SLAVE19_WUSER    = SLAVE_WUSER[(19+1)*USER_WIDTH-1:19*USER_WIDTH];  
      assign  SLAVE19_WVALID   = SLAVE_WVALID[19];      
      assign  SLAVE19_BREADY   = SLAVE_BREADY[19];        
      assign  SLAVE19_ARID     = SLAVE_ARID[(19+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:19*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE19_ARADDR   = SLAVE_ARADDR[(19+1)*ADDR_WIDTH-1:19*ADDR_WIDTH];  
      assign  SLAVE19_ARLEN    = SLAVE_ARLEN[(19+1)*8-1:19*8];  
      assign  SLAVE19_ARSIZE   = SLAVE_ARSIZE[(19+1)*3-1:19*3];  
      assign  SLAVE19_ARBURST  = SLAVE_ARBURST[(19+1)*2-1:19*2];  
      assign  SLAVE19_ARLOCK   = SLAVE_ARLOCK[(19+1)*2-1:19*2];  
      assign  SLAVE19_ARCACHE  = SLAVE_ARCACHE[(19+1)*4-1:19*4] ;  
      assign  SLAVE19_ARPROT   = SLAVE_ARPROT[(19+1)*3-1:19*3] ;  
      assign  SLAVE19_ARREGION = SLAVE_ARREGION[(19+1)*4-1:19*4];   
      assign  SLAVE19_ARQOS    = SLAVE_ARQOS[(19+1)*4-1:19*4];  
      assign  SLAVE19_ARUSER   = SLAVE_ARUSER[(19+1)*USER_WIDTH-1:19*USER_WIDTH];  
      assign  SLAVE19_ARVALID  = SLAVE_ARVALID[19];      
      assign  SLAVE19_RREADY   = SLAVE_RREADY[19];  

      //Inputs      
      assign  SLAVE_AWREADY[19]                                                                    = SLAVE19_AWREADY;          
      assign  SLAVE_WREADY[19]                                                                     = SLAVE19_WREADY;        
      assign  SLAVE_BID[(19+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:19*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE19_BID;  
      assign  SLAVE_BRESP[(19+1)*2-1:19*2]                                                         = SLAVE19_BRESP;  
      assign  SLAVE_BUSER[(19+1)*USER_WIDTH-1:19*USER_WIDTH]                                       = SLAVE19_BUSER;  
      assign  SLAVE_BVALID[19]                                                                     = SLAVE19_BVALID;        
      assign  SLAVE_ARREADY[19]                                                                    = SLAVE19_ARREADY;        
      assign  SLAVE_RID[(19+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:19*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE19_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(19+1)*13-1:13*19]-1:SDW_LOWER_VEC[(19+1)*13-1:13*19]]     = SLAVE19_RDATA;  
      assign  SLAVE_RRESP[(19+1)*2-1:19*2]                                                         = SLAVE19_RRESP;  
      assign  SLAVE_RLAST[19]                                                                      = SLAVE19_RLAST;  
      assign  SLAVE_RUSER[(19+1)*USER_WIDTH-1:19*USER_WIDTH]                                       = SLAVE19_RUSER;  
      assign  SLAVE_RVALID[19]                                                                     = SLAVE19_RVALID;
    end
    
    if ( NUM_SLAVES > 20 )
    begin
      //===================================================================
      //Slave20 Combine Signals
      //===================================================================
      //======================= SLAVE20 TO/FROM External Side=================
      //Outputs
      assign  SLAVE20_AWID     = SLAVE_AWID[(20+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:20*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE20_AWADDR   = SLAVE_AWADDR[(20+1)*ADDR_WIDTH-1:20*ADDR_WIDTH];  
      assign  SLAVE20_AWLEN    = SLAVE_AWLEN[(20+1)*8-1:20*8];  
      assign  SLAVE20_AWSIZE   = SLAVE_AWSIZE[(20+1)*3-1:20*3];  
      assign  SLAVE20_AWBURST  = SLAVE_AWBURST[(20+1)*2-1:20*2];  
      assign  SLAVE20_AWLOCK   = SLAVE_AWLOCK[(20+1)*2-1:20*2];  
      assign  SLAVE20_AWCACHE  = SLAVE_AWCACHE[(20+1)*4-1:20*4];  
      assign  SLAVE20_AWPROT   = SLAVE_AWPROT[(20+1)*3-1:20*3];  
      assign  SLAVE20_AWREGION = SLAVE_AWREGION[(20+1)*4-1:20*4];   
      assign  SLAVE20_AWQOS    = SLAVE_AWQOS[(20+1)*4-1:20*4];  
      assign  SLAVE20_AWUSER   = SLAVE_AWUSER[(20+1)*USER_WIDTH-1:20*USER_WIDTH];  
      assign  SLAVE20_AWVALID  = SLAVE_AWVALID[20];  
      assign  SLAVE20_WID      = SLAVE_WID[(20+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:20*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE20_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(20+1)*13-1:13*20]-1:SDW_LOWER_VEC[(20+1)*13-1:13*20]];  
      assign  SLAVE20_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(20+1)*13-1:13*20]/8-1:SDW_LOWER_VEC[(20+1)*13-1:13*20]/8];  
      assign  SLAVE20_WLAST    = SLAVE_WLAST[20];  
      assign  SLAVE20_WUSER    = SLAVE_WUSER[(20+1)*USER_WIDTH-1:20*USER_WIDTH];  
      assign  SLAVE20_WVALID   = SLAVE_WVALID[20];      
      assign  SLAVE20_BREADY   = SLAVE_BREADY[20];        
      assign  SLAVE20_ARID     = SLAVE_ARID[(20+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:20*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE20_ARADDR   = SLAVE_ARADDR[(20+1)*ADDR_WIDTH-1:20*ADDR_WIDTH];  
      assign  SLAVE20_ARLEN    = SLAVE_ARLEN[(20+1)*8-1:20*8];  
      assign  SLAVE20_ARSIZE   = SLAVE_ARSIZE[(20+1)*3-1:20*3];  
      assign  SLAVE20_ARBURST  = SLAVE_ARBURST[(20+1)*2-1:20*2];  
      assign  SLAVE20_ARLOCK   = SLAVE_ARLOCK[(20+1)*2-1:20*2];  
      assign  SLAVE20_ARCACHE  = SLAVE_ARCACHE[(20+1)*4-1:20*4] ;  
      assign  SLAVE20_ARPROT   = SLAVE_ARPROT[(20+1)*3-1:20*3] ;  
      assign  SLAVE20_ARREGION = SLAVE_ARREGION[(20+1)*4-1:20*4];   
      assign  SLAVE20_ARQOS    = SLAVE_ARQOS[(20+1)*4-1:20*4];  
      assign  SLAVE20_ARUSER   = SLAVE_ARUSER[(20+1)*USER_WIDTH-1:20*USER_WIDTH];  
      assign  SLAVE20_ARVALID  = SLAVE_ARVALID[20];      
      assign  SLAVE20_RREADY   = SLAVE_RREADY[20];  

      //Inputs      
      assign  SLAVE_AWREADY[20]                                                                    = SLAVE20_AWREADY;          
      assign  SLAVE_WREADY[20]                                                                     = SLAVE20_WREADY;        
      assign  SLAVE_BID[(20+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:20*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE20_BID;  
      assign  SLAVE_BRESP[(20+1)*2-1:20*2]                                                         = SLAVE20_BRESP;  
      assign  SLAVE_BUSER[(20+1)*USER_WIDTH-1:20*USER_WIDTH]                                       = SLAVE20_BUSER;  
      assign  SLAVE_BVALID[20]                                                                     = SLAVE20_BVALID;        
      assign  SLAVE_ARREADY[20]                                                                    = SLAVE20_ARREADY;        
      assign  SLAVE_RID[(20+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:20*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE20_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(20+1)*13-1:13*20]-1:SDW_LOWER_VEC[(20+1)*13-1:13*20]]     = SLAVE20_RDATA;  
      assign  SLAVE_RRESP[(20+1)*2-1:20*2]                                                         = SLAVE20_RRESP;  
      assign  SLAVE_RLAST[20]                                                                      = SLAVE20_RLAST;  
      assign  SLAVE_RUSER[(20+1)*USER_WIDTH-1:20*USER_WIDTH]                                       = SLAVE20_RUSER;  
      assign  SLAVE_RVALID[20]                                                                     = SLAVE20_RVALID;
    end
    
    if ( NUM_SLAVES > 21 )
    begin
      //===================================================================
      //Slave21 Combine Signals
      //===================================================================
      //======================= SLAVE21 TO/FROM External Side=================
      //Outputs
      assign  SLAVE21_AWID     = SLAVE_AWID[(21+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:21*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE21_AWADDR   = SLAVE_AWADDR[(21+1)*ADDR_WIDTH-1:21*ADDR_WIDTH];  
      assign  SLAVE21_AWLEN    = SLAVE_AWLEN[(21+1)*8-1:21*8];  
      assign  SLAVE21_AWSIZE   = SLAVE_AWSIZE[(21+1)*3-1:21*3];  
      assign  SLAVE21_AWBURST  = SLAVE_AWBURST[(21+1)*2-1:21*2];  
      assign  SLAVE21_AWLOCK   = SLAVE_AWLOCK[(21+1)*2-1:21*2];  
      assign  SLAVE21_AWCACHE  = SLAVE_AWCACHE[(21+1)*4-1:21*4];  
      assign  SLAVE21_AWPROT   = SLAVE_AWPROT[(21+1)*3-1:21*3];  
      assign  SLAVE21_AWREGION = SLAVE_AWREGION[(21+1)*4-1:21*4];   
      assign  SLAVE21_AWQOS    = SLAVE_AWQOS[(21+1)*4-1:21*4];  
      assign  SLAVE21_AWUSER   = SLAVE_AWUSER[(21+1)*USER_WIDTH-1:21*USER_WIDTH];  
      assign  SLAVE21_AWVALID  = SLAVE_AWVALID[21];  
      assign  SLAVE21_WID      = SLAVE_WID[(21+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:21*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE21_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(21+1)*13-1:13*21]-1:SDW_LOWER_VEC[(21+1)*13-1:13*21]];  
      assign  SLAVE21_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(21+1)*13-1:13*21]/8-1:SDW_LOWER_VEC[(21+1)*13-1:13*21]/8];  
      assign  SLAVE21_WLAST    = SLAVE_WLAST[21];  
      assign  SLAVE21_WUSER    = SLAVE_WUSER[(21+1)*USER_WIDTH-1:21*USER_WIDTH];  
      assign  SLAVE21_WVALID   = SLAVE_WVALID[21];      
      assign  SLAVE21_BREADY   = SLAVE_BREADY[21];        
      assign  SLAVE21_ARID     = SLAVE_ARID[(21+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:21*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE21_ARADDR   = SLAVE_ARADDR[(21+1)*ADDR_WIDTH-1:21*ADDR_WIDTH];  
      assign  SLAVE21_ARLEN    = SLAVE_ARLEN[(21+1)*8-1:21*8];  
      assign  SLAVE21_ARSIZE   = SLAVE_ARSIZE[(21+1)*3-1:21*3];  
      assign  SLAVE21_ARBURST  = SLAVE_ARBURST[(21+1)*2-1:21*2];  
      assign  SLAVE21_ARLOCK   = SLAVE_ARLOCK[(21+1)*2-1:21*2];  
      assign  SLAVE21_ARCACHE  = SLAVE_ARCACHE[(21+1)*4-1:21*4] ;  
      assign  SLAVE21_ARPROT   = SLAVE_ARPROT[(21+1)*3-1:21*3] ;  
      assign  SLAVE21_ARREGION = SLAVE_ARREGION[(21+1)*4-1:21*4];   
      assign  SLAVE21_ARQOS    = SLAVE_ARQOS[(21+1)*4-1:21*4];  
      assign  SLAVE21_ARUSER   = SLAVE_ARUSER[(21+1)*USER_WIDTH-1:21*USER_WIDTH];  
      assign  SLAVE21_ARVALID  = SLAVE_ARVALID[21];      
      assign  SLAVE21_RREADY   = SLAVE_RREADY[21];  

      //Inputs      
      assign  SLAVE_AWREADY[21]                                                                    = SLAVE21_AWREADY;          
      assign  SLAVE_WREADY[21]                                                                     = SLAVE21_WREADY;        
      assign  SLAVE_BID[(21+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:21*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE21_BID;  
      assign  SLAVE_BRESP[(21+1)*2-1:21*2]                                                         = SLAVE21_BRESP;  
      assign  SLAVE_BUSER[(21+1)*USER_WIDTH-1:21*USER_WIDTH]                                       = SLAVE21_BUSER;  
      assign  SLAVE_BVALID[21]                                                                     = SLAVE21_BVALID;        
      assign  SLAVE_ARREADY[21]                                                                    = SLAVE21_ARREADY;        
      assign  SLAVE_RID[(21+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:21*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE21_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(21+1)*13-1:13*21]-1:SDW_LOWER_VEC[(21+1)*13-1:13*21]]     = SLAVE21_RDATA;  
      assign  SLAVE_RRESP[(21+1)*2-1:21*2]                                                         = SLAVE21_RRESP;  
      assign  SLAVE_RLAST[21]                                                                      = SLAVE21_RLAST;  
      assign  SLAVE_RUSER[(21+1)*USER_WIDTH-1:21*USER_WIDTH]                                       = SLAVE21_RUSER;  
      assign  SLAVE_RVALID[21]                                                                     = SLAVE21_RVALID;
    end
    
    if ( NUM_SLAVES > 22 )
    begin
      //===================================================================
      //Slave22 Combine Signals
      //===================================================================
      //======================= SLAVE22 TO/FROM External Side=================
      //Outputs
      assign  SLAVE22_AWID     = SLAVE_AWID[(22+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:22*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE22_AWADDR   = SLAVE_AWADDR[(22+1)*ADDR_WIDTH-1:22*ADDR_WIDTH];  
      assign  SLAVE22_AWLEN    = SLAVE_AWLEN[(22+1)*8-1:22*8];  
      assign  SLAVE22_AWSIZE   = SLAVE_AWSIZE[(22+1)*3-1:22*3];  
      assign  SLAVE22_AWBURST  = SLAVE_AWBURST[(22+1)*2-1:22*2];  
      assign  SLAVE22_AWLOCK   = SLAVE_AWLOCK[(22+1)*2-1:22*2];  
      assign  SLAVE22_AWCACHE  = SLAVE_AWCACHE[(22+1)*4-1:22*4];  
      assign  SLAVE22_AWPROT   = SLAVE_AWPROT[(22+1)*3-1:22*3];  
      assign  SLAVE22_AWREGION = SLAVE_AWREGION[(22+1)*4-1:22*4];   
      assign  SLAVE22_AWQOS    = SLAVE_AWQOS[(22+1)*4-1:22*4];  
      assign  SLAVE22_AWUSER   = SLAVE_AWUSER[(22+1)*USER_WIDTH-1:22*USER_WIDTH];  
      assign  SLAVE22_AWVALID  = SLAVE_AWVALID[22];  
      assign  SLAVE22_WID      = SLAVE_WID[(22+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:22*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE22_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(22+1)*13-1:13*22]-1:SDW_LOWER_VEC[(22+1)*13-1:13*22]];  
      assign  SLAVE22_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(22+1)*13-1:13*22]/8-1:SDW_LOWER_VEC[(22+1)*13-1:13*22]/8];  
      assign  SLAVE22_WLAST    = SLAVE_WLAST[22];  
      assign  SLAVE22_WUSER    = SLAVE_WUSER[(22+1)*USER_WIDTH-1:22*USER_WIDTH];  
      assign  SLAVE22_WVALID   = SLAVE_WVALID[22];      
      assign  SLAVE22_BREADY   = SLAVE_BREADY[22];        
      assign  SLAVE22_ARID     = SLAVE_ARID[(22+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:22*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE22_ARADDR   = SLAVE_ARADDR[(22+1)*ADDR_WIDTH-1:22*ADDR_WIDTH];  
      assign  SLAVE22_ARLEN    = SLAVE_ARLEN[(22+1)*8-1:22*8];  
      assign  SLAVE22_ARSIZE   = SLAVE_ARSIZE[(22+1)*3-1:22*3];  
      assign  SLAVE22_ARBURST  = SLAVE_ARBURST[(22+1)*2-1:22*2];  
      assign  SLAVE22_ARLOCK   = SLAVE_ARLOCK[(22+1)*2-1:22*2];  
      assign  SLAVE22_ARCACHE  = SLAVE_ARCACHE[(22+1)*4-1:22*4] ;  
      assign  SLAVE22_ARPROT   = SLAVE_ARPROT[(22+1)*3-1:22*3] ;  
      assign  SLAVE22_ARREGION = SLAVE_ARREGION[(22+1)*4-1:22*4];   
      assign  SLAVE22_ARQOS    = SLAVE_ARQOS[(22+1)*4-1:22*4];  
      assign  SLAVE22_ARUSER   = SLAVE_ARUSER[(22+1)*USER_WIDTH-1:22*USER_WIDTH];  
      assign  SLAVE22_ARVALID  = SLAVE_ARVALID[22];      
      assign  SLAVE22_RREADY   = SLAVE_RREADY[22];  

      //Inputs      
      assign  SLAVE_AWREADY[22]                                                                    = SLAVE22_AWREADY;          
      assign  SLAVE_WREADY[22]                                                                     = SLAVE22_WREADY;        
      assign  SLAVE_BID[(22+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:22*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE22_BID;  
      assign  SLAVE_BRESP[(22+1)*2-1:22*2]                                                         = SLAVE22_BRESP;  
      assign  SLAVE_BUSER[(22+1)*USER_WIDTH-1:22*USER_WIDTH]                                       = SLAVE22_BUSER;  
      assign  SLAVE_BVALID[22]                                                                     = SLAVE22_BVALID;        
      assign  SLAVE_ARREADY[22]                                                                    = SLAVE22_ARREADY;        
      assign  SLAVE_RID[(22+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:22*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE22_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(22+1)*13-1:13*22]-1:SDW_LOWER_VEC[(22+1)*13-1:13*22]]     = SLAVE22_RDATA;  
      assign  SLAVE_RRESP[(22+1)*2-1:22*2]                                                         = SLAVE22_RRESP;  
      assign  SLAVE_RLAST[22]                                                                      = SLAVE22_RLAST;  
      assign  SLAVE_RUSER[(22+1)*USER_WIDTH-1:22*USER_WIDTH]                                       = SLAVE22_RUSER;  
      assign  SLAVE_RVALID[22]                                                                     = SLAVE22_RVALID;
    end
    
    if ( NUM_SLAVES > 23 )
    begin
      //===================================================================
      //Slave23 Combine Signals
      //===================================================================
      //======================= SLAVE23 TO/FROM External Side=================
      //Outputs
      assign  SLAVE23_AWID     = SLAVE_AWID[(23+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:23*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE23_AWADDR   = SLAVE_AWADDR[(23+1)*ADDR_WIDTH-1:23*ADDR_WIDTH];  
      assign  SLAVE23_AWLEN    = SLAVE_AWLEN[(23+1)*8-1:23*8];  
      assign  SLAVE23_AWSIZE   = SLAVE_AWSIZE[(23+1)*3-1:23*3];  
      assign  SLAVE23_AWBURST  = SLAVE_AWBURST[(23+1)*2-1:23*2];  
      assign  SLAVE23_AWLOCK   = SLAVE_AWLOCK[(23+1)*2-1:23*2];  
      assign  SLAVE23_AWCACHE  = SLAVE_AWCACHE[(23+1)*4-1:23*4];  
      assign  SLAVE23_AWPROT   = SLAVE_AWPROT[(23+1)*3-1:23*3];  
      assign  SLAVE23_AWREGION = SLAVE_AWREGION[(23+1)*4-1:23*4];   
      assign  SLAVE23_AWQOS    = SLAVE_AWQOS[(23+1)*4-1:23*4];  
      assign  SLAVE23_AWUSER   = SLAVE_AWUSER[(23+1)*USER_WIDTH-1:23*USER_WIDTH];  
      assign  SLAVE23_AWVALID  = SLAVE_AWVALID[23];  
      assign  SLAVE23_WID      = SLAVE_WID[(23+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:23*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE23_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(23+1)*13-1:13*23]-1:SDW_LOWER_VEC[(23+1)*13-1:13*23]];  
      assign  SLAVE23_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(23+1)*13-1:13*23]/8-1:SDW_LOWER_VEC[(23+1)*13-1:13*23]/8];  
      assign  SLAVE23_WLAST    = SLAVE_WLAST[23];  
      assign  SLAVE23_WUSER    = SLAVE_WUSER[(23+1)*USER_WIDTH-1:23*USER_WIDTH];  
      assign  SLAVE23_WVALID   = SLAVE_WVALID[23];      
      assign  SLAVE23_BREADY   = SLAVE_BREADY[23];        
      assign  SLAVE23_ARID     = SLAVE_ARID[(23+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:23*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE23_ARADDR   = SLAVE_ARADDR[(23+1)*ADDR_WIDTH-1:23*ADDR_WIDTH];  
      assign  SLAVE23_ARLEN    = SLAVE_ARLEN[(23+1)*8-1:23*8];  
      assign  SLAVE23_ARSIZE   = SLAVE_ARSIZE[(23+1)*3-1:23*3];  
      assign  SLAVE23_ARBURST  = SLAVE_ARBURST[(23+1)*2-1:23*2];  
      assign  SLAVE23_ARLOCK   = SLAVE_ARLOCK[(23+1)*2-1:23*2];  
      assign  SLAVE23_ARCACHE  = SLAVE_ARCACHE[(23+1)*4-1:23*4] ;  
      assign  SLAVE23_ARPROT   = SLAVE_ARPROT[(23+1)*3-1:23*3] ;  
      assign  SLAVE23_ARREGION = SLAVE_ARREGION[(23+1)*4-1:23*4];   
      assign  SLAVE23_ARQOS    = SLAVE_ARQOS[(23+1)*4-1:23*4];  
      assign  SLAVE23_ARUSER   = SLAVE_ARUSER[(23+1)*USER_WIDTH-1:23*USER_WIDTH];  
      assign  SLAVE23_ARVALID  = SLAVE_ARVALID[23];      
      assign  SLAVE23_RREADY   = SLAVE_RREADY[23];  

      //Inputs      
      assign  SLAVE_AWREADY[23]                                                                    = SLAVE23_AWREADY;          
      assign  SLAVE_WREADY[23]                                                                     = SLAVE23_WREADY;        
      assign  SLAVE_BID[(23+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:23*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE23_BID;  
      assign  SLAVE_BRESP[(23+1)*2-1:23*2]                                                         = SLAVE23_BRESP;  
      assign  SLAVE_BUSER[(23+1)*USER_WIDTH-1:23*USER_WIDTH]                                       = SLAVE23_BUSER;  
      assign  SLAVE_BVALID[23]                                                                     = SLAVE23_BVALID;        
      assign  SLAVE_ARREADY[23]                                                                    = SLAVE23_ARREADY;        
      assign  SLAVE_RID[(23+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:23*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE23_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(23+1)*13-1:13*23]-1:SDW_LOWER_VEC[(23+1)*13-1:13*23]]     = SLAVE23_RDATA;  
      assign  SLAVE_RRESP[(23+1)*2-1:23*2]                                                         = SLAVE23_RRESP;  
      assign  SLAVE_RLAST[23]                                                                      = SLAVE23_RLAST;  
      assign  SLAVE_RUSER[(23+1)*USER_WIDTH-1:23*USER_WIDTH]                                       = SLAVE23_RUSER;  
      assign  SLAVE_RVALID[23]                                                                     = SLAVE23_RVALID;
    end
    
    if ( NUM_SLAVES > 24 )
    begin
      //===================================================================
      //Slave24 Combine Signals
      //===================================================================
      //======================= SLAVE24 TO/FROM External Side=================
      //Outputs
      assign  SLAVE24_AWID     = SLAVE_AWID[(24+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:24*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE24_AWADDR   = SLAVE_AWADDR[(24+1)*ADDR_WIDTH-1:24*ADDR_WIDTH];  
      assign  SLAVE24_AWLEN    = SLAVE_AWLEN[(24+1)*8-1:24*8];  
      assign  SLAVE24_AWSIZE   = SLAVE_AWSIZE[(24+1)*3-1:24*3];  
      assign  SLAVE24_AWBURST  = SLAVE_AWBURST[(24+1)*2-1:24*2];  
      assign  SLAVE24_AWLOCK   = SLAVE_AWLOCK[(24+1)*2-1:24*2];  
      assign  SLAVE24_AWCACHE  = SLAVE_AWCACHE[(24+1)*4-1:24*4];  
      assign  SLAVE24_AWPROT   = SLAVE_AWPROT[(24+1)*3-1:24*3];  
      assign  SLAVE24_AWREGION = SLAVE_AWREGION[(24+1)*4-1:24*4];   
      assign  SLAVE24_AWQOS    = SLAVE_AWQOS[(24+1)*4-1:24*4];  
      assign  SLAVE24_AWUSER   = SLAVE_AWUSER[(24+1)*USER_WIDTH-1:24*USER_WIDTH];  
      assign  SLAVE24_AWVALID  = SLAVE_AWVALID[24];  
      assign  SLAVE24_WID      = SLAVE_WID[(24+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:24*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE24_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(24+1)*13-1:13*24]-1:SDW_LOWER_VEC[(24+1)*13-1:13*24]];  
      assign  SLAVE24_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(24+1)*13-1:13*24]/8-1:SDW_LOWER_VEC[(24+1)*13-1:13*24]/8];  
      assign  SLAVE24_WLAST    = SLAVE_WLAST[24];  
      assign  SLAVE24_WUSER    = SLAVE_WUSER[(24+1)*USER_WIDTH-1:24*USER_WIDTH];  
      assign  SLAVE24_WVALID   = SLAVE_WVALID[24];      
      assign  SLAVE24_BREADY   = SLAVE_BREADY[24];        
      assign  SLAVE24_ARID     = SLAVE_ARID[(24+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:24*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE24_ARADDR   = SLAVE_ARADDR[(24+1)*ADDR_WIDTH-1:24*ADDR_WIDTH];  
      assign  SLAVE24_ARLEN    = SLAVE_ARLEN[(24+1)*8-1:24*8];  
      assign  SLAVE24_ARSIZE   = SLAVE_ARSIZE[(24+1)*3-1:24*3];  
      assign  SLAVE24_ARBURST  = SLAVE_ARBURST[(24+1)*2-1:24*2];  
      assign  SLAVE24_ARLOCK   = SLAVE_ARLOCK[(24+1)*2-1:24*2];  
      assign  SLAVE24_ARCACHE  = SLAVE_ARCACHE[(24+1)*4-1:24*4] ;  
      assign  SLAVE24_ARPROT   = SLAVE_ARPROT[(24+1)*3-1:24*3] ;  
      assign  SLAVE24_ARREGION = SLAVE_ARREGION[(24+1)*4-1:24*4];   
      assign  SLAVE24_ARQOS    = SLAVE_ARQOS[(24+1)*4-1:24*4];  
      assign  SLAVE24_ARUSER   = SLAVE_ARUSER[(24+1)*USER_WIDTH-1:24*USER_WIDTH];  
      assign  SLAVE24_ARVALID  = SLAVE_ARVALID[24];      
      assign  SLAVE24_RREADY   = SLAVE_RREADY[24];  

      //Inputs      
      assign  SLAVE_AWREADY[24]                                                                    = SLAVE24_AWREADY;          
      assign  SLAVE_WREADY[24]                                                                     = SLAVE24_WREADY;        
      assign  SLAVE_BID[(24+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:24*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE24_BID;  
      assign  SLAVE_BRESP[(24+1)*2-1:24*2]                                                         = SLAVE24_BRESP;  
      assign  SLAVE_BUSER[(24+1)*USER_WIDTH-1:24*USER_WIDTH]                                       = SLAVE24_BUSER;  
      assign  SLAVE_BVALID[24]                                                                     = SLAVE24_BVALID;        
      assign  SLAVE_ARREADY[24]                                                                    = SLAVE24_ARREADY;        
      assign  SLAVE_RID[(24+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:24*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE24_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(24+1)*13-1:13*24]-1:SDW_LOWER_VEC[(24+1)*13-1:13*24]]     = SLAVE24_RDATA;  
      assign  SLAVE_RRESP[(24+1)*2-1:24*2]                                                         = SLAVE24_RRESP;  
      assign  SLAVE_RLAST[24]                                                                      = SLAVE24_RLAST;  
      assign  SLAVE_RUSER[(24+1)*USER_WIDTH-1:24*USER_WIDTH]                                       = SLAVE24_RUSER;  
      assign  SLAVE_RVALID[24]                                                                     = SLAVE24_RVALID;
    end
    
    if ( NUM_SLAVES > 25 )
    begin
      //===================================================================
      //Slave25 Combine Signals
      //===================================================================
      //======================= SLAVE25 TO/FROM External Side=================
      //Outputs
      assign  SLAVE25_AWID     = SLAVE_AWID[(25+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:25*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE25_AWADDR   = SLAVE_AWADDR[(25+1)*ADDR_WIDTH-1:25*ADDR_WIDTH];  
      assign  SLAVE25_AWLEN    = SLAVE_AWLEN[(25+1)*8-1:25*8];  
      assign  SLAVE25_AWSIZE   = SLAVE_AWSIZE[(25+1)*3-1:25*3];  
      assign  SLAVE25_AWBURST  = SLAVE_AWBURST[(25+1)*2-1:25*2];  
      assign  SLAVE25_AWLOCK   = SLAVE_AWLOCK[(25+1)*2-1:25*2];  
      assign  SLAVE25_AWCACHE  = SLAVE_AWCACHE[(25+1)*4-1:25*4];  
      assign  SLAVE25_AWPROT   = SLAVE_AWPROT[(25+1)*3-1:25*3];  
      assign  SLAVE25_AWREGION = SLAVE_AWREGION[(25+1)*4-1:25*4];   
      assign  SLAVE25_AWQOS    = SLAVE_AWQOS[(25+1)*4-1:25*4];  
      assign  SLAVE25_AWUSER   = SLAVE_AWUSER[(25+1)*USER_WIDTH-1:25*USER_WIDTH];  
      assign  SLAVE25_AWVALID  = SLAVE_AWVALID[25];  
      assign  SLAVE25_WID      = SLAVE_WID[(25+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:25*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE25_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(25+1)*13-1:13*25]-1:SDW_LOWER_VEC[(25+1)*13-1:13*25]];  
      assign  SLAVE25_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(25+1)*13-1:13*25]/8-1:SDW_LOWER_VEC[(25+1)*13-1:13*25]/8];  
      assign  SLAVE25_WLAST    = SLAVE_WLAST[25];  
      assign  SLAVE25_WUSER    = SLAVE_WUSER[(25+1)*USER_WIDTH-1:25*USER_WIDTH];  
      assign  SLAVE25_WVALID   = SLAVE_WVALID[25];      
      assign  SLAVE25_BREADY   = SLAVE_BREADY[25];        
      assign  SLAVE25_ARID     = SLAVE_ARID[(25+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:25*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE25_ARADDR   = SLAVE_ARADDR[(25+1)*ADDR_WIDTH-1:25*ADDR_WIDTH];  
      assign  SLAVE25_ARLEN    = SLAVE_ARLEN[(25+1)*8-1:25*8];  
      assign  SLAVE25_ARSIZE   = SLAVE_ARSIZE[(25+1)*3-1:25*3];  
      assign  SLAVE25_ARBURST  = SLAVE_ARBURST[(25+1)*2-1:25*2];  
      assign  SLAVE25_ARLOCK   = SLAVE_ARLOCK[(25+1)*2-1:25*2];  
      assign  SLAVE25_ARCACHE  = SLAVE_ARCACHE[(25+1)*4-1:25*4] ;  
      assign  SLAVE25_ARPROT   = SLAVE_ARPROT[(25+1)*3-1:25*3] ;  
      assign  SLAVE25_ARREGION = SLAVE_ARREGION[(25+1)*4-1:25*4];   
      assign  SLAVE25_ARQOS    = SLAVE_ARQOS[(25+1)*4-1:25*4];  
      assign  SLAVE25_ARUSER   = SLAVE_ARUSER[(25+1)*USER_WIDTH-1:25*USER_WIDTH];  
      assign  SLAVE25_ARVALID  = SLAVE_ARVALID[25];      
      assign  SLAVE25_RREADY   = SLAVE_RREADY[25];  

      //Inputs      
      assign  SLAVE_AWREADY[25]                                                                    = SLAVE25_AWREADY;          
      assign  SLAVE_WREADY[25]                                                                     = SLAVE25_WREADY;        
      assign  SLAVE_BID[(25+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:25*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE25_BID;  
      assign  SLAVE_BRESP[(25+1)*2-1:25*2]                                                         = SLAVE25_BRESP;  
      assign  SLAVE_BUSER[(25+1)*USER_WIDTH-1:25*USER_WIDTH]                                       = SLAVE25_BUSER;  
      assign  SLAVE_BVALID[25]                                                                     = SLAVE25_BVALID;        
      assign  SLAVE_ARREADY[25]                                                                    = SLAVE25_ARREADY;        
      assign  SLAVE_RID[(25+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:25*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE25_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(25+1)*13-1:13*25]-1:SDW_LOWER_VEC[(25+1)*13-1:13*25]]     = SLAVE25_RDATA;  
      assign  SLAVE_RRESP[(25+1)*2-1:25*2]                                                         = SLAVE25_RRESP;  
      assign  SLAVE_RLAST[25]                                                                      = SLAVE25_RLAST;  
      assign  SLAVE_RUSER[(25+1)*USER_WIDTH-1:25*USER_WIDTH]                                       = SLAVE25_RUSER;  
      assign  SLAVE_RVALID[25]                                                                     = SLAVE25_RVALID;
    end
    
    if ( NUM_SLAVES > 26 )
    begin
      //===================================================================
      //Slave26 Combine Signals
      //===================================================================
      //======================= SLAVE26 TO/FROM External Side=================
      //Outputs
      assign  SLAVE26_AWID     = SLAVE_AWID[(26+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:26*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE26_AWADDR   = SLAVE_AWADDR[(26+1)*ADDR_WIDTH-1:26*ADDR_WIDTH];  
      assign  SLAVE26_AWLEN    = SLAVE_AWLEN[(26+1)*8-1:26*8];  
      assign  SLAVE26_AWSIZE   = SLAVE_AWSIZE[(26+1)*3-1:26*3];  
      assign  SLAVE26_AWBURST  = SLAVE_AWBURST[(26+1)*2-1:26*2];  
      assign  SLAVE26_AWLOCK   = SLAVE_AWLOCK[(26+1)*2-1:26*2];  
      assign  SLAVE26_AWCACHE  = SLAVE_AWCACHE[(26+1)*4-1:26*4];  
      assign  SLAVE26_AWPROT   = SLAVE_AWPROT[(26+1)*3-1:26*3];  
      assign  SLAVE26_AWREGION = SLAVE_AWREGION[(26+1)*4-1:26*4];   
      assign  SLAVE26_AWQOS    = SLAVE_AWQOS[(26+1)*4-1:26*4];  
      assign  SLAVE26_AWUSER   = SLAVE_AWUSER[(26+1)*USER_WIDTH-1:26*USER_WIDTH];  
      assign  SLAVE26_AWVALID  = SLAVE_AWVALID[26];  
      assign  SLAVE26_WID      = SLAVE_WID[(26+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:26*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE26_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(26+1)*13-1:13*26]-1:SDW_LOWER_VEC[(26+1)*13-1:13*26]];  
      assign  SLAVE26_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(26+1)*13-1:13*26]/8-1:SDW_LOWER_VEC[(26+1)*13-1:13*26]/8];  
      assign  SLAVE26_WLAST    = SLAVE_WLAST[26];  
      assign  SLAVE26_WUSER    = SLAVE_WUSER[(26+1)*USER_WIDTH-1:26*USER_WIDTH];  
      assign  SLAVE26_WVALID   = SLAVE_WVALID[26];      
      assign  SLAVE26_BREADY   = SLAVE_BREADY[26];        
      assign  SLAVE26_ARID     = SLAVE_ARID[(26+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:26*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE26_ARADDR   = SLAVE_ARADDR[(26+1)*ADDR_WIDTH-1:26*ADDR_WIDTH];  
      assign  SLAVE26_ARLEN    = SLAVE_ARLEN[(26+1)*8-1:26*8];  
      assign  SLAVE26_ARSIZE   = SLAVE_ARSIZE[(26+1)*3-1:26*3];  
      assign  SLAVE26_ARBURST  = SLAVE_ARBURST[(26+1)*2-1:26*2];  
      assign  SLAVE26_ARLOCK   = SLAVE_ARLOCK[(26+1)*2-1:26*2];  
      assign  SLAVE26_ARCACHE  = SLAVE_ARCACHE[(26+1)*4-1:26*4] ;  
      assign  SLAVE26_ARPROT   = SLAVE_ARPROT[(26+1)*3-1:26*3] ;  
      assign  SLAVE26_ARREGION = SLAVE_ARREGION[(26+1)*4-1:26*4];   
      assign  SLAVE26_ARQOS    = SLAVE_ARQOS[(26+1)*4-1:26*4];  
      assign  SLAVE26_ARUSER   = SLAVE_ARUSER[(26+1)*USER_WIDTH-1:26*USER_WIDTH];  
      assign  SLAVE26_ARVALID  = SLAVE_ARVALID[26];      
      assign  SLAVE26_RREADY   = SLAVE_RREADY[26];  

      //Inputs      
      assign  SLAVE_AWREADY[26]                                                                    = SLAVE26_AWREADY;          
      assign  SLAVE_WREADY[26]                                                                     = SLAVE26_WREADY;        
      assign  SLAVE_BID[(26+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:26*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE26_BID;  
      assign  SLAVE_BRESP[(26+1)*2-1:26*2]                                                         = SLAVE26_BRESP;  
      assign  SLAVE_BUSER[(26+1)*USER_WIDTH-1:26*USER_WIDTH]                                       = SLAVE26_BUSER;  
      assign  SLAVE_BVALID[26]                                                                     = SLAVE26_BVALID;        
      assign  SLAVE_ARREADY[26]                                                                    = SLAVE26_ARREADY;        
      assign  SLAVE_RID[(26+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:26*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE26_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(26+1)*13-1:13*26]-1:SDW_LOWER_VEC[(26+1)*13-1:13*26]]     = SLAVE26_RDATA;  
      assign  SLAVE_RRESP[(26+1)*2-1:26*2]                                                         = SLAVE26_RRESP;  
      assign  SLAVE_RLAST[26]                                                                      = SLAVE26_RLAST;  
      assign  SLAVE_RUSER[(26+1)*USER_WIDTH-1:26*USER_WIDTH]                                       = SLAVE26_RUSER;  
      assign  SLAVE_RVALID[26]                                                                     = SLAVE26_RVALID;
    end
    
    if ( NUM_SLAVES > 27 )
    begin
      //===================================================================
      //Slave27 Combine Signals
      //===================================================================
      //======================= SLAVE27 TO/FROM External Side=================
      //Outputs
      assign  SLAVE27_AWID     = SLAVE_AWID[(27+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:27*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE27_AWADDR   = SLAVE_AWADDR[(27+1)*ADDR_WIDTH-1:27*ADDR_WIDTH];  
      assign  SLAVE27_AWLEN    = SLAVE_AWLEN[(27+1)*8-1:27*8];  
      assign  SLAVE27_AWSIZE   = SLAVE_AWSIZE[(27+1)*3-1:27*3];  
      assign  SLAVE27_AWBURST  = SLAVE_AWBURST[(27+1)*2-1:27*2];  
      assign  SLAVE27_AWLOCK   = SLAVE_AWLOCK[(27+1)*2-1:27*2];  
      assign  SLAVE27_AWCACHE  = SLAVE_AWCACHE[(27+1)*4-1:27*4];  
      assign  SLAVE27_AWPROT   = SLAVE_AWPROT[(27+1)*3-1:27*3];  
      assign  SLAVE27_AWREGION = SLAVE_AWREGION[(27+1)*4-1:27*4];   
      assign  SLAVE27_AWQOS    = SLAVE_AWQOS[(27+1)*4-1:27*4];  
      assign  SLAVE27_AWUSER   = SLAVE_AWUSER[(27+1)*USER_WIDTH-1:27*USER_WIDTH];  
      assign  SLAVE27_AWVALID  = SLAVE_AWVALID[27];  
      assign  SLAVE27_WID      = SLAVE_WID[(27+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:27*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE27_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(27+1)*13-1:13*27]-1:SDW_LOWER_VEC[(27+1)*13-1:13*27]];  
      assign  SLAVE27_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(27+1)*13-1:13*27]/8-1:SDW_LOWER_VEC[(27+1)*13-1:13*27]/8];  
      assign  SLAVE27_WLAST    = SLAVE_WLAST[27];  
      assign  SLAVE27_WUSER    = SLAVE_WUSER[(27+1)*USER_WIDTH-1:27*USER_WIDTH];  
      assign  SLAVE27_WVALID   = SLAVE_WVALID[27];      
      assign  SLAVE27_BREADY   = SLAVE_BREADY[27];        
      assign  SLAVE27_ARID     = SLAVE_ARID[(27+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:27*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE27_ARADDR   = SLAVE_ARADDR[(27+1)*ADDR_WIDTH-1:27*ADDR_WIDTH];  
      assign  SLAVE27_ARLEN    = SLAVE_ARLEN[(27+1)*8-1:27*8];  
      assign  SLAVE27_ARSIZE   = SLAVE_ARSIZE[(27+1)*3-1:27*3];  
      assign  SLAVE27_ARBURST  = SLAVE_ARBURST[(27+1)*2-1:27*2];  
      assign  SLAVE27_ARLOCK   = SLAVE_ARLOCK[(27+1)*2-1:27*2];  
      assign  SLAVE27_ARCACHE  = SLAVE_ARCACHE[(27+1)*4-1:27*4] ;  
      assign  SLAVE27_ARPROT   = SLAVE_ARPROT[(27+1)*3-1:27*3] ;  
      assign  SLAVE27_ARREGION = SLAVE_ARREGION[(27+1)*4-1:27*4];   
      assign  SLAVE27_ARQOS    = SLAVE_ARQOS[(27+1)*4-1:27*4];  
      assign  SLAVE27_ARUSER   = SLAVE_ARUSER[(27+1)*USER_WIDTH-1:27*USER_WIDTH];  
      assign  SLAVE27_ARVALID  = SLAVE_ARVALID[27];      
      assign  SLAVE27_RREADY   = SLAVE_RREADY[27];  

      //Inputs      
      assign  SLAVE_AWREADY[27]                                                                    = SLAVE27_AWREADY;          
      assign  SLAVE_WREADY[27]                                                                     = SLAVE27_WREADY;        
      assign  SLAVE_BID[(27+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:27*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE27_BID;  
      assign  SLAVE_BRESP[(27+1)*2-1:27*2]                                                         = SLAVE27_BRESP;  
      assign  SLAVE_BUSER[(27+1)*USER_WIDTH-1:27*USER_WIDTH]                                       = SLAVE27_BUSER;  
      assign  SLAVE_BVALID[27]                                                                     = SLAVE27_BVALID;        
      assign  SLAVE_ARREADY[27]                                                                    = SLAVE27_ARREADY;        
      assign  SLAVE_RID[(27+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:27*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE27_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(27+1)*13-1:13*27]-1:SDW_LOWER_VEC[(27+1)*13-1:13*27]]     = SLAVE27_RDATA;  
      assign  SLAVE_RRESP[(27+1)*2-1:27*2]                                                         = SLAVE27_RRESP;  
      assign  SLAVE_RLAST[27]                                                                      = SLAVE27_RLAST;  
      assign  SLAVE_RUSER[(27+1)*USER_WIDTH-1:27*USER_WIDTH]                                       = SLAVE27_RUSER;  
      assign  SLAVE_RVALID[27]                                                                     = SLAVE27_RVALID;
    end
    
    if ( NUM_SLAVES > 28 )
    begin
      //===================================================================
      //Slave28 Combine Signals
      //===================================================================
      //======================= SLAVE28 TO/FROM External Side=================
      //Outputs
      assign  SLAVE28_AWID     = SLAVE_AWID[(28+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:28*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE28_AWADDR   = SLAVE_AWADDR[(28+1)*ADDR_WIDTH-1:28*ADDR_WIDTH];  
      assign  SLAVE28_AWLEN    = SLAVE_AWLEN[(28+1)*8-1:28*8];  
      assign  SLAVE28_AWSIZE   = SLAVE_AWSIZE[(28+1)*3-1:28*3];  
      assign  SLAVE28_AWBURST  = SLAVE_AWBURST[(28+1)*2-1:28*2];  
      assign  SLAVE28_AWLOCK   = SLAVE_AWLOCK[(28+1)*2-1:28*2];  
      assign  SLAVE28_AWCACHE  = SLAVE_AWCACHE[(28+1)*4-1:28*4];  
      assign  SLAVE28_AWPROT   = SLAVE_AWPROT[(28+1)*3-1:28*3];  
      assign  SLAVE28_AWREGION = SLAVE_AWREGION[(28+1)*4-1:28*4];   
      assign  SLAVE28_AWQOS    = SLAVE_AWQOS[(28+1)*4-1:28*4];  
      assign  SLAVE28_AWUSER   = SLAVE_AWUSER[(28+1)*USER_WIDTH-1:28*USER_WIDTH];  
      assign  SLAVE28_AWVALID  = SLAVE_AWVALID[28];  
      assign  SLAVE28_WID      = SLAVE_WID[(28+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:28*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE28_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(28+1)*13-1:13*28]-1:SDW_LOWER_VEC[(28+1)*13-1:13*28]];  
      assign  SLAVE28_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(28+1)*13-1:13*28]/8-1:SDW_LOWER_VEC[(28+1)*13-1:13*28]/8];  
      assign  SLAVE28_WLAST    = SLAVE_WLAST[28];  
      assign  SLAVE28_WUSER    = SLAVE_WUSER[(28+1)*USER_WIDTH-1:28*USER_WIDTH];  
      assign  SLAVE28_WVALID   = SLAVE_WVALID[28];      
      assign  SLAVE28_BREADY   = SLAVE_BREADY[28];        
      assign  SLAVE28_ARID     = SLAVE_ARID[(28+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:28*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE28_ARADDR   = SLAVE_ARADDR[(28+1)*ADDR_WIDTH-1:28*ADDR_WIDTH];  
      assign  SLAVE28_ARLEN    = SLAVE_ARLEN[(28+1)*8-1:28*8];  
      assign  SLAVE28_ARSIZE   = SLAVE_ARSIZE[(28+1)*3-1:28*3];  
      assign  SLAVE28_ARBURST  = SLAVE_ARBURST[(28+1)*2-1:28*2];  
      assign  SLAVE28_ARLOCK   = SLAVE_ARLOCK[(28+1)*2-1:28*2];  
      assign  SLAVE28_ARCACHE  = SLAVE_ARCACHE[(28+1)*4-1:28*4] ;  
      assign  SLAVE28_ARPROT   = SLAVE_ARPROT[(28+1)*3-1:28*3] ;  
      assign  SLAVE28_ARREGION = SLAVE_ARREGION[(28+1)*4-1:28*4];   
      assign  SLAVE28_ARQOS    = SLAVE_ARQOS[(28+1)*4-1:28*4];  
      assign  SLAVE28_ARUSER   = SLAVE_ARUSER[(28+1)*USER_WIDTH-1:28*USER_WIDTH];  
      assign  SLAVE28_ARVALID  = SLAVE_ARVALID[28];      
      assign  SLAVE28_RREADY   = SLAVE_RREADY[28];  

      //Inputs      
      assign  SLAVE_AWREADY[28]                                                                    = SLAVE28_AWREADY;          
      assign  SLAVE_WREADY[28]                                                                     = SLAVE28_WREADY;        
      assign  SLAVE_BID[(28+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:28*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE28_BID;  
      assign  SLAVE_BRESP[(28+1)*2-1:28*2]                                                         = SLAVE28_BRESP;  
      assign  SLAVE_BUSER[(28+1)*USER_WIDTH-1:28*USER_WIDTH]                                       = SLAVE28_BUSER;  
      assign  SLAVE_BVALID[28]                                                                     = SLAVE28_BVALID;        
      assign  SLAVE_ARREADY[28]                                                                    = SLAVE28_ARREADY;        
      assign  SLAVE_RID[(28+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:28*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE28_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(28+1)*13-1:13*28]-1:SDW_LOWER_VEC[(28+1)*13-1:13*28]]     = SLAVE28_RDATA;  
      assign  SLAVE_RRESP[(28+1)*2-1:28*2]                                                         = SLAVE28_RRESP;  
      assign  SLAVE_RLAST[28]                                                                      = SLAVE28_RLAST;  
      assign  SLAVE_RUSER[(28+1)*USER_WIDTH-1:28*USER_WIDTH]                                       = SLAVE28_RUSER;  
      assign  SLAVE_RVALID[28]                                                                     = SLAVE28_RVALID;
    end
    
    if ( NUM_SLAVES > 29 )
    begin
      //===================================================================
      //Slave29 Combine Signals
      //===================================================================
      //======================= SLAVE29 TO/FROM External Side=================
      //Outputs
      assign  SLAVE29_AWID     = SLAVE_AWID[(29+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:29*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE29_AWADDR   = SLAVE_AWADDR[(29+1)*ADDR_WIDTH-1:29*ADDR_WIDTH];  
      assign  SLAVE29_AWLEN    = SLAVE_AWLEN[(29+1)*8-1:29*8];  
      assign  SLAVE29_AWSIZE   = SLAVE_AWSIZE[(29+1)*3-1:29*3];  
      assign  SLAVE29_AWBURST  = SLAVE_AWBURST[(29+1)*2-1:29*2];  
      assign  SLAVE29_AWLOCK   = SLAVE_AWLOCK[(29+1)*2-1:29*2];  
      assign  SLAVE29_AWCACHE  = SLAVE_AWCACHE[(29+1)*4-1:29*4];  
      assign  SLAVE29_AWPROT   = SLAVE_AWPROT[(29+1)*3-1:29*3];  
      assign  SLAVE29_AWREGION = SLAVE_AWREGION[(29+1)*4-1:29*4];   
      assign  SLAVE29_AWQOS    = SLAVE_AWQOS[(29+1)*4-1:29*4];  
      assign  SLAVE29_AWUSER   = SLAVE_AWUSER[(29+1)*USER_WIDTH-1:29*USER_WIDTH];  
      assign  SLAVE29_AWVALID  = SLAVE_AWVALID[29];  
      assign  SLAVE29_WID      = SLAVE_WID[(29+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:29*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE29_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(29+1)*13-1:13*29]-1:SDW_LOWER_VEC[(29+1)*13-1:13*29]];  
      assign  SLAVE29_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(29+1)*13-1:13*29]/8-1:SDW_LOWER_VEC[(29+1)*13-1:13*29]/8];  
      assign  SLAVE29_WLAST    = SLAVE_WLAST[29];  
      assign  SLAVE29_WUSER    = SLAVE_WUSER[(29+1)*USER_WIDTH-1:29*USER_WIDTH];  
      assign  SLAVE29_WVALID   = SLAVE_WVALID[29];      
      assign  SLAVE29_BREADY   = SLAVE_BREADY[29];        
      assign  SLAVE29_ARID     = SLAVE_ARID[(29+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:29*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE29_ARADDR   = SLAVE_ARADDR[(29+1)*ADDR_WIDTH-1:29*ADDR_WIDTH];  
      assign  SLAVE29_ARLEN    = SLAVE_ARLEN[(29+1)*8-1:29*8];  
      assign  SLAVE29_ARSIZE   = SLAVE_ARSIZE[(29+1)*3-1:29*3];  
      assign  SLAVE29_ARBURST  = SLAVE_ARBURST[(29+1)*2-1:29*2];  
      assign  SLAVE29_ARLOCK   = SLAVE_ARLOCK[(29+1)*2-1:29*2];  
      assign  SLAVE29_ARCACHE  = SLAVE_ARCACHE[(29+1)*4-1:29*4] ;  
      assign  SLAVE29_ARPROT   = SLAVE_ARPROT[(29+1)*3-1:29*3] ;  
      assign  SLAVE29_ARREGION = SLAVE_ARREGION[(29+1)*4-1:29*4];   
      assign  SLAVE29_ARQOS    = SLAVE_ARQOS[(29+1)*4-1:29*4];  
      assign  SLAVE29_ARUSER   = SLAVE_ARUSER[(29+1)*USER_WIDTH-1:29*USER_WIDTH];  
      assign  SLAVE29_ARVALID  = SLAVE_ARVALID[29];      
      assign  SLAVE29_RREADY   = SLAVE_RREADY[29];  

      //Inputs      
      assign  SLAVE_AWREADY[29]                                                                    = SLAVE29_AWREADY;          
      assign  SLAVE_WREADY[29]                                                                     = SLAVE29_WREADY;        
      assign  SLAVE_BID[(29+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:29*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE29_BID;  
      assign  SLAVE_BRESP[(29+1)*2-1:29*2]                                                         = SLAVE29_BRESP;  
      assign  SLAVE_BUSER[(29+1)*USER_WIDTH-1:29*USER_WIDTH]                                       = SLAVE29_BUSER;  
      assign  SLAVE_BVALID[29]                                                                     = SLAVE29_BVALID;        
      assign  SLAVE_ARREADY[29]                                                                    = SLAVE29_ARREADY;        
      assign  SLAVE_RID[(29+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:29*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE29_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(29+1)*13-1:13*29]-1:SDW_LOWER_VEC[(29+1)*13-1:13*29]]     = SLAVE29_RDATA;  
      assign  SLAVE_RRESP[(29+1)*2-1:29*2]                                                         = SLAVE29_RRESP;  
      assign  SLAVE_RLAST[29]                                                                      = SLAVE29_RLAST;  
      assign  SLAVE_RUSER[(29+1)*USER_WIDTH-1:29*USER_WIDTH]                                       = SLAVE29_RUSER;  
      assign  SLAVE_RVALID[29]                                                                     = SLAVE29_RVALID;
    end
    
    if ( NUM_SLAVES > 30 )
    begin
      //===================================================================
      //Slave30 Combine Signals
      //===================================================================
      //======================= SLAVE30 TO/FROM External Side=================
      //Outputs
      assign  SLAVE30_AWID     = SLAVE_AWID[(30+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:30*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE30_AWADDR   = SLAVE_AWADDR[(30+1)*ADDR_WIDTH-1:30*ADDR_WIDTH];  
      assign  SLAVE30_AWLEN    = SLAVE_AWLEN[(30+1)*8-1:30*8];  
      assign  SLAVE30_AWSIZE   = SLAVE_AWSIZE[(30+1)*3-1:30*3];  
      assign  SLAVE30_AWBURST  = SLAVE_AWBURST[(30+1)*2-1:30*2];  
      assign  SLAVE30_AWLOCK   = SLAVE_AWLOCK[(30+1)*2-1:30*2];  
      assign  SLAVE30_AWCACHE  = SLAVE_AWCACHE[(30+1)*4-1:30*4];  
      assign  SLAVE30_AWPROT   = SLAVE_AWPROT[(30+1)*3-1:30*3];  
      assign  SLAVE30_AWREGION = SLAVE_AWREGION[(30+1)*4-1:30*4];   
      assign  SLAVE30_AWQOS    = SLAVE_AWQOS[(30+1)*4-1:30*4];  
      assign  SLAVE30_AWUSER   = SLAVE_AWUSER[(30+1)*USER_WIDTH-1:30*USER_WIDTH];  
      assign  SLAVE30_AWVALID  = SLAVE_AWVALID[30];  
      assign  SLAVE30_WID      = SLAVE_WID[(30+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:30*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE30_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(30+1)*13-1:13*30]-1:SDW_LOWER_VEC[(30+1)*13-1:13*30]];  
      assign  SLAVE30_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(30+1)*13-1:13*30]/8-1:SDW_LOWER_VEC[(30+1)*13-1:13*30]/8];  
      assign  SLAVE30_WLAST    = SLAVE_WLAST[30];  
      assign  SLAVE30_WUSER    = SLAVE_WUSER[(30+1)*USER_WIDTH-1:30*USER_WIDTH];  
      assign  SLAVE30_WVALID   = SLAVE_WVALID[30];      
      assign  SLAVE30_BREADY   = SLAVE_BREADY[30];        
      assign  SLAVE30_ARID     = SLAVE_ARID[(30+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:30*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE30_ARADDR   = SLAVE_ARADDR[(30+1)*ADDR_WIDTH-1:30*ADDR_WIDTH];  
      assign  SLAVE30_ARLEN    = SLAVE_ARLEN[(30+1)*8-1:30*8];  
      assign  SLAVE30_ARSIZE   = SLAVE_ARSIZE[(30+1)*3-1:30*3];  
      assign  SLAVE30_ARBURST  = SLAVE_ARBURST[(30+1)*2-1:30*2];  
      assign  SLAVE30_ARLOCK   = SLAVE_ARLOCK[(30+1)*2-1:30*2];  
      assign  SLAVE30_ARCACHE  = SLAVE_ARCACHE[(30+1)*4-1:30*4] ;  
      assign  SLAVE30_ARPROT   = SLAVE_ARPROT[(30+1)*3-1:30*3] ;  
      assign  SLAVE30_ARREGION = SLAVE_ARREGION[(30+1)*4-1:30*4];   
      assign  SLAVE30_ARQOS    = SLAVE_ARQOS[(30+1)*4-1:30*4];  
      assign  SLAVE30_ARUSER   = SLAVE_ARUSER[(30+1)*USER_WIDTH-1:30*USER_WIDTH];  
      assign  SLAVE30_ARVALID  = SLAVE_ARVALID[30];      
      assign  SLAVE30_RREADY   = SLAVE_RREADY[30];  

      //Inputs      
      assign  SLAVE_AWREADY[30]                                                                    = SLAVE30_AWREADY;          
      assign  SLAVE_WREADY[30]                                                                     = SLAVE30_WREADY;        
      assign  SLAVE_BID[(30+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:30*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE30_BID;  
      assign  SLAVE_BRESP[(30+1)*2-1:30*2]                                                         = SLAVE30_BRESP;  
      assign  SLAVE_BUSER[(30+1)*USER_WIDTH-1:30*USER_WIDTH]                                       = SLAVE30_BUSER;  
      assign  SLAVE_BVALID[30]                                                                     = SLAVE30_BVALID;        
      assign  SLAVE_ARREADY[30]                                                                    = SLAVE30_ARREADY;        
      assign  SLAVE_RID[(30+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:30*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE30_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(30+1)*13-1:13*30]-1:SDW_LOWER_VEC[(30+1)*13-1:13*30]]     = SLAVE30_RDATA;  
      assign  SLAVE_RRESP[(30+1)*2-1:30*2]                                                         = SLAVE30_RRESP;  
      assign  SLAVE_RLAST[30]                                                                      = SLAVE30_RLAST;  
      assign  SLAVE_RUSER[(30+1)*USER_WIDTH-1:30*USER_WIDTH]                                       = SLAVE30_RUSER;  
      assign  SLAVE_RVALID[30]                                                                     = SLAVE30_RVALID;
    end
    
    if ( NUM_SLAVES > 31 )
    begin
      //===================================================================
      //Slave31 Combine Signals
      //===================================================================
      //======================= SLAVE31 TO/FROM External Side=================
      //Outputs
      assign  SLAVE31_AWID     = SLAVE_AWID[(31+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:31*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE31_AWADDR   = SLAVE_AWADDR[(31+1)*ADDR_WIDTH-1:31*ADDR_WIDTH];  
      assign  SLAVE31_AWLEN    = SLAVE_AWLEN[(31+1)*8-1:31*8];  
      assign  SLAVE31_AWSIZE   = SLAVE_AWSIZE[(31+1)*3-1:31*3];  
      assign  SLAVE31_AWBURST  = SLAVE_AWBURST[(31+1)*2-1:31*2];  
      assign  SLAVE31_AWLOCK   = SLAVE_AWLOCK[(31+1)*2-1:31*2];  
      assign  SLAVE31_AWCACHE  = SLAVE_AWCACHE[(31+1)*4-1:31*4];  
      assign  SLAVE31_AWPROT   = SLAVE_AWPROT[(31+1)*3-1:31*3];  
      assign  SLAVE31_AWREGION = SLAVE_AWREGION[(31+1)*4-1:31*4];   
      assign  SLAVE31_AWQOS    = SLAVE_AWQOS[(31+1)*4-1:31*4];  
      assign  SLAVE31_AWUSER   = SLAVE_AWUSER[(31+1)*USER_WIDTH-1:31*USER_WIDTH];  
      assign  SLAVE31_AWVALID  = SLAVE_AWVALID[31];  
      assign  SLAVE31_WID      = SLAVE_WID[(31+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:31*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE31_WDATA    = SLAVE_WDATA[SDW_UPPER_VEC[(31+1)*13-1:13*31]-1:SDW_LOWER_VEC[(31+1)*13-1:13*31]];  
      assign  SLAVE31_WSTRB    = SLAVE_WSTRB[SDW_UPPER_VEC[(31+1)*13-1:13*31]/8-1:SDW_LOWER_VEC[(31+1)*13-1:13*31]/8];  
      assign  SLAVE31_WLAST    = SLAVE_WLAST[31];  
      assign  SLAVE31_WUSER    = SLAVE_WUSER[(31+1)*USER_WIDTH-1:31*USER_WIDTH];  
      assign  SLAVE31_WVALID   = SLAVE_WVALID[31];      
      assign  SLAVE31_BREADY   = SLAVE_BREADY[31];        
      assign  SLAVE31_ARID     = SLAVE_ARID[(31+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:31*(NUM_MASTERS_WIDTH+ID_WIDTH)];  
      assign  SLAVE31_ARADDR   = SLAVE_ARADDR[(31+1)*ADDR_WIDTH-1:31*ADDR_WIDTH];  
      assign  SLAVE31_ARLEN    = SLAVE_ARLEN[(31+1)*8-1:31*8];  
      assign  SLAVE31_ARSIZE   = SLAVE_ARSIZE[(31+1)*3-1:31*3];  
      assign  SLAVE31_ARBURST  = SLAVE_ARBURST[(31+1)*2-1:31*2];  
      assign  SLAVE31_ARLOCK   = SLAVE_ARLOCK[(31+1)*2-1:31*2];  
      assign  SLAVE31_ARCACHE  = SLAVE_ARCACHE[(31+1)*4-1:31*4] ;  
      assign  SLAVE31_ARPROT   = SLAVE_ARPROT[(31+1)*3-1:31*3] ;  
      assign  SLAVE31_ARREGION = SLAVE_ARREGION[(31+1)*4-1:31*4];   
      assign  SLAVE31_ARQOS    = SLAVE_ARQOS[(31+1)*4-1:31*4];  
      assign  SLAVE31_ARUSER   = SLAVE_ARUSER[(31+1)*USER_WIDTH-1:31*USER_WIDTH];  
      assign  SLAVE31_ARVALID  = SLAVE_ARVALID[31];      
      assign  SLAVE31_RREADY   = SLAVE_RREADY[31];  

      //Inputs      
      assign  SLAVE_AWREADY[31]                                                                    = SLAVE31_AWREADY;          
      assign  SLAVE_WREADY[31]                                                                     = SLAVE31_WREADY;        
      assign  SLAVE_BID[(31+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:31*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE31_BID;  
      assign  SLAVE_BRESP[(31+1)*2-1:31*2]                                                         = SLAVE31_BRESP;  
      assign  SLAVE_BUSER[(31+1)*USER_WIDTH-1:31*USER_WIDTH]                                       = SLAVE31_BUSER;  
      assign  SLAVE_BVALID[31]                                                                     = SLAVE31_BVALID;        
      assign  SLAVE_ARREADY[31]                                                                    = SLAVE31_ARREADY;        
      assign  SLAVE_RID[(31+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:31*(NUM_MASTERS_WIDTH+ID_WIDTH)]     = SLAVE31_RID;  
      assign  SLAVE_RDATA[SDW_UPPER_VEC[(31+1)*13-1:13*31]-1:SDW_LOWER_VEC[(31+1)*13-1:13*31]]     = SLAVE31_RDATA;  
      assign  SLAVE_RRESP[(31+1)*2-1:31*2]                                                         = SLAVE31_RRESP;  
      assign  SLAVE_RLAST[31]                                                                      = SLAVE31_RLAST;  
      assign  SLAVE_RUSER[(31+1)*USER_WIDTH-1:31*USER_WIDTH]                                       = SLAVE31_RUSER;  
      assign  SLAVE_RVALID[31]                                                                     = SLAVE31_RVALID;
    end
    
  //===============================================================================================================================

  // Master clocks
  generate
  if(MASTER0_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[0] = M_CLK0;
  else
    assign M_CLK[0] = ACLK;
  endgenerate
  
  generate
  if(MASTER1_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[1] = M_CLK1;
  else
    assign M_CLK[1] = ACLK;
  endgenerate
  
  generate
  if(MASTER2_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[2] = M_CLK2;
  else
    assign M_CLK[2] = ACLK;
  endgenerate
  
  generate
  if(MASTER3_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[3] = M_CLK3;
  else
    assign M_CLK[3] = ACLK;
  endgenerate
  
  generate
  if(MASTER4_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[4] = M_CLK4;
  else
    assign M_CLK[4] = ACLK;
  endgenerate
  
  generate
  if(MASTER5_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[5] = M_CLK5;
  else
    assign M_CLK[5] = ACLK;
  endgenerate
  
  generate
  if(MASTER6_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[6] = M_CLK6;
  else
    assign M_CLK[6] = ACLK;
  endgenerate
  
  generate
  if(MASTER7_CLOCK_DOMAIN_CROSSING)
    assign M_CLK[7] = M_CLK7;
  else
    assign M_CLK[7] = ACLK;
  endgenerate
  
  // Slave Clocks
  generate
  if(SLAVE0_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[0] = S_CLK0;
  else
    assign S_CLK[0] = ACLK;
  endgenerate
  
  generate
  if(SLAVE1_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[1] = S_CLK1;
  else
    assign S_CLK[1] = ACLK;
  endgenerate
  
  generate
  if(SLAVE2_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[2] = S_CLK2;
  else
    assign S_CLK[2] = ACLK;
  endgenerate
  
  generate
  if(SLAVE3_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[3] = S_CLK3;
  else
    assign S_CLK[3] = ACLK;
  endgenerate
  
  generate
  if(SLAVE4_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[4] = S_CLK4;
  else
    assign S_CLK[4] = ACLK;
  endgenerate
  
  generate
  if(SLAVE5_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[5] = S_CLK5;
  else
    assign S_CLK[5] = ACLK;
  endgenerate
  
  generate
  if(SLAVE6_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[6] = S_CLK6;
  else
    assign S_CLK[6] = ACLK;
  endgenerate
  
  generate
  if(SLAVE7_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[7] = S_CLK7;
  else
    assign S_CLK[7] = ACLK;
  endgenerate
  
  generate
  if(SLAVE8_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[8] = S_CLK8;
  else
    assign S_CLK[8] = ACLK;
  endgenerate
  
  generate
  if(SLAVE9_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[9] = S_CLK9;
  else
    assign S_CLK[9] = ACLK;
  endgenerate
  
  generate
  if(SLAVE10_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[10] = S_CLK10;
  else
    assign S_CLK[10] = ACLK;
  endgenerate

  generate
  if(SLAVE11_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[11] = S_CLK11;
  else
    assign S_CLK[11] = ACLK;
  endgenerate

  generate
  if(SLAVE12_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[12] = S_CLK12;
  else
    assign S_CLK[12] = ACLK;
  endgenerate
  
  generate
  if(SLAVE13_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[13] = S_CLK13;
  else
    assign S_CLK[13] = ACLK;
  endgenerate

  generate
  if(SLAVE14_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[14] = S_CLK14;
  else
    assign S_CLK[14] = ACLK;
  endgenerate
  
  generate
  if(SLAVE15_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[15] = S_CLK15;
  else
    assign S_CLK[15] = ACLK;
  endgenerate

  generate
  if(SLAVE16_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[16] = S_CLK16;
  else
    assign S_CLK[16] = ACLK;
  endgenerate

  generate
  if(SLAVE17_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[17] = S_CLK17;
  else
    assign S_CLK[17] = ACLK;
  endgenerate

  generate
  if(SLAVE18_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[18] = S_CLK18;
  else
    assign S_CLK[18] = ACLK;
  endgenerate

  generate
  if(SLAVE19_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[19] = S_CLK19;
  else
    assign S_CLK[19] = ACLK;
  endgenerate

  generate
  if(SLAVE20_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[20] = S_CLK20;
  else
    assign S_CLK[20] = ACLK;
  endgenerate

  generate
  if(SLAVE21_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[21] = S_CLK21;
  else
    assign S_CLK[21] = ACLK;
  endgenerate

  generate
  if(SLAVE22_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[22] = S_CLK22;
  else
    assign S_CLK[22] = ACLK;
  endgenerate

  generate
  if(SLAVE23_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[23] = S_CLK23;
  else
    assign S_CLK[23] = ACLK;
  endgenerate

  generate
  if(SLAVE24_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[24] = S_CLK24;
  else
    assign S_CLK[24] = ACLK;
  endgenerate

  generate
  if(SLAVE25_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[25] = S_CLK25;
  else
    assign S_CLK[25] = ACLK;
  endgenerate

  generate
  if(SLAVE26_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[26] = S_CLK26;
  else
    assign S_CLK[26] = ACLK;
  endgenerate

  generate
  if(SLAVE27_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[27] = S_CLK27;
  else
    assign S_CLK[27] = ACLK;
  endgenerate

  generate
  if(SLAVE28_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[28] = S_CLK28;
  else
    assign S_CLK[28] = ACLK;
  endgenerate

  generate
  if(SLAVE29_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[29] = S_CLK29;
  else
    assign S_CLK[29] = ACLK;
  endgenerate

  generate
  if(SLAVE30_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[30] = S_CLK30;
  else
    assign S_CLK[30] = ACLK;
  endgenerate

  generate
  if(SLAVE31_CLOCK_DOMAIN_CROSSING)
    assign S_CLK[31] = S_CLK31;
  else
    assign S_CLK[31] = ACLK;
  endgenerate

  //Reset synchronizer to remove cdc violations
  
  caxi4interconnect_ResetSycnc arst_aclk_sync
  (
    .sysClk	( ACLK ),
	.sysReset_L( ARESETN ),			// active low reset synchronoise to RE AClk - asserted async.
	.sysReset( ACLK_syncReset  )	// active low sysReset synchronised to ACLK
  );
  
  caxi4interconnect_Axi4CrossBar #
    (
      .FAMILY                      (  19  ), 
      .NUM_MASTERS                 ( NUM_MASTERS ),         // defines number of masters
      .NUM_MASTERS_WIDTH           ( NUM_MASTERS_WIDTH ),
      .NUM_SLAVES                  ( NUM_SLAVES ),         // defines number of slaves

      .ADDR_WIDTH                  ( ADDR_WIDTH  ),        
      .DATA_WIDTH                  ( DATA_WIDTH  ),
      .ID_WIDTH                    ( ID_WIDTH ),

      .NUM_THREADS                 ( NUM_THREADS ),
      .OPEN_TRANS_MAX              ( OPEN_TRANS_MAX ), 
      .OPEN_WRTRANS_MAX            ( OPEN_WRTRANS_MAX ),
      .OPEN_RDTRANS_MAX            ( OPEN_RDTRANS_MAX ),

      .UPPER_COMPARE_BIT           ( UPPER_COMPARE_BIT ),
      .LOWER_COMPARE_BIT           ( LOWER_COMPARE_BIT ),

      .SLOT_BASE_VEC               ( SLOT_BASE_VEC ),
      .SLOT_MIN_VEC                ( SLOT_MIN_VEC ),
      .SLOT_MAX_VEC                ( SLOT_MAX_VEC ),
    
      .SUPPORT_USER_SIGNALS        ( SUPPORT_USER_SIGNALS ),
      .USER_WIDTH                  ( USER_WIDTH ),
      .CROSSBAR_MODE               ( CROSSBAR_MODE ),

      .MASTER_WRITE_CONNECTIVITY   ( MASTER_WRITE_CONNECTIVITY ), 
      .MASTER_READ_CONNECTIVITY    ( MASTER_READ_CONNECTIVITY  ),
      .HI_FREQ                     ( HI_FREQ ),
      .RD_ARB_EN                   ( RD_ARB_EN )
    )
  axicb (
      // Global Signals
      .ACLK    ( ACLK ),
      .ARESETN ( ACLK_syncReset ),
  
      // Master Write Address Ports
      .MASTER_AWID     ( masterAWID ),
      .MASTER_AWADDR   ( masterAWADDR ),
      .MASTER_AWLEN    ( masterAWLEN ),
      .MASTER_AWSIZE   ( masterAWSIZE ),
      .MASTER_AWBURST  ( masterAWBURST ),
      .MASTER_AWLOCK   ( masterAWLOCK ),
      .MASTER_AWCACHE  ( masterAWCACHE ),
      .MASTER_AWPROT   ( masterAWPROT ),
      .MASTER_AWREGION ( masterAWREGION ),
      .MASTER_AWQOS    ( masterAWQOS ),        // not used
      .MASTER_AWUSER   ( masterAWUSER ),        // not used
      .MASTER_AWVALID  ( masterAWVALID ),
      .MASTER_AWREADY  ( masterAWREADY ),

      // Master Write Data Ports
      .MASTER_WDATA   ( masterWDATA ),
      .MASTER_WSTRB   ( masterWSTRB ),
      .MASTER_WLAST   ( masterWLAST ),
      .MASTER_WUSER   ( masterWUSER ),
      .MASTER_WVALID  ( masterWVALID ),
      .MASTER_WREADY  ( masterWREADY ),
 
      // Master Write Response Ports
      .MASTER_BID     ( masterBID ),
      .MASTER_BRESP   ( masterBRESP ),
      .MASTER_BUSER   ( masterBUSER ),
      .MASTER_BVALID  ( masterBVALID ),
      .MASTER_BREADY  ( masterBREADY ),

      // Master Read Address Ports
      .MASTER_ARID     ( masterARID ),
      .MASTER_ARADDR   ( masterARADDR ),
      .MASTER_ARLEN    ( masterARLEN ),
      .MASTER_ARSIZE   ( masterARSIZE ),
      .MASTER_ARBURST  ( masterARBURST ),
      .MASTER_ARLOCK   ( masterARLOCK ),
      .MASTER_ARCACHE  ( masterARCACHE ),
      .MASTER_ARPROT   ( masterARPROT ),
      .MASTER_ARREGION ( masterARREGION ),
      .MASTER_ARQOS    ( masterARQOS ),        // not used
      .MASTER_ARUSER   ( masterARUSER ),
      .MASTER_ARVALID  ( masterARVALID ),
      .MASTER_ARREADY  ( masterARREADY ),

      // Master Read Data Ports
      .MASTER_RID     ( masterRID ),
      .MASTER_RDATA   ( masterRDATA ), // output from this module, masterRDATA = slaveRDATA
      .MASTER_RRESP   ( masterRRESP ),
      .MASTER_RLAST   ( masterRLAST ),
      .MASTER_RUSER   ( masterRUSER ),
      .MASTER_RVALID  ( masterRVALID ),
      .MASTER_RREADY  ( masterRREADY ),
   
      // Slave Write Address Port
      .SLAVE_AWID      ( slaveAWID ),
      .SLAVE_AWADDR    ( slaveAWADDR ),
      .SLAVE_AWLEN     ( slaveAWLEN ),
      .SLAVE_AWSIZE    ( slaveAWSIZE ),
      .SLAVE_AWBURST   ( slaveAWBURST ),
      .SLAVE_AWLOCK    ( slaveAWLOCK ),
      .SLAVE_AWCACHE   ( slaveAWCACHE ),
      .SLAVE_AWPROT    ( slaveAWPROT ),
      .SLAVE_AWREGION  ( slaveAWREGION ),      // not used
      .SLAVE_AWQOS     ( slaveAWQOS ),      // not used
      .SLAVE_AWUSER    ( slaveAWUSER ),
      .SLAVE_AWVALID   ( slaveAWVALID ),
      .SLAVE_AWREADY   ( slaveAWREADY ),
   
      // Slave Write Data Ports
      .SLAVE_WDATA   ( slaveWDATA ),
      .SLAVE_WSTRB   ( slaveWSTRB ),
      .SLAVE_WLAST   ( slaveWLAST ),
      .SLAVE_WUSER   ( slaveWUSER ),
      .SLAVE_WVALID  ( slaveWVALID ),
      .SLAVE_WREADY  ( slaveWREADY ),

      // Slave Write Response Ports
      .SLAVE_BID     ( slaveBID ),
      .SLAVE_BRESP   ( slaveBRESP ),
      .SLAVE_BUSER   ( slaveBUSER ),
      .SLAVE_BVALID  ( slaveBVALID ),
      .SLAVE_BREADY  ( slaveBREADY ),
   
      // Slave Read Address Port
      .SLAVE_ARID      ( slaveARID ),
      .SLAVE_ARADDR    ( slaveARADDR ),
      .SLAVE_ARLEN     ( slaveARLEN ),
      .SLAVE_ARSIZE    ( slaveARSIZE ),
      .SLAVE_ARBURST   ( slaveARBURST ),
      .SLAVE_ARLOCK    ( slaveARLOCK ),
      .SLAVE_ARCACHE   ( slaveARCACHE ),
      .SLAVE_ARPROT    ( slaveARPROT ),
      .SLAVE_ARREGION  ( slaveARREGION ),      // not used
      .SLAVE_ARQOS     ( slaveARQOS ),      // not used
      .SLAVE_ARUSER    ( slaveARUSER ),
      .SLAVE_ARVALID   ( slaveARVALID ),
      .SLAVE_ARREADY   ( slaveARREADY ),
   
      // Slave Read Data Ports
      .SLAVE_RID     ( slaveRID ),
      .SLAVE_RDATA   ( slaveRDATA ), // input to this module
      .SLAVE_RRESP   ( slaveRRESP ),
      .SLAVE_RLAST   ( slaveRLAST ),
      .SLAVE_RUSER   ( slaveRUSER ),      // not used
      .SLAVE_RVALID  ( slaveRVALID ),
      .SLAVE_RREADY  ( slaveRREADY )
   );
   
  //===============================================================================================================================
        genvar mst;
  generate
                for (mst=0; mst<NUM_MASTERS; mst=mst+1) begin : MstConvertor_loop
    caxi4interconnect_MasterConvertor #
          (
            .DEF_BURST_LEN          ( MASTER_DEF_BURST_LEN[(mst+1)*8-1:mst*8] ),
            .DWC_DATA_FIFO_DEPTH    ( MASTER_DWC_DATA_FIFO_DEPTH[(mst+1)*14-1:mst*14] ),
            .DWC_ADDR_FIFO_DEPTH_CEILING (DWC_ADDR_FIFO_DEPTH_CEILING),
            .MASTER_TYPE            ( MASTER_TYPE [(mst+1)*2-1:mst*2] ) ,   // Protocol type = AXI4 - 2'b00, AXI4Lite - 2'b01, AXI3 - 2'b10
            .MASTER_NUMBER          ( mst ),          // master number
            .AWCHAN_RS              ( MASTER_AWCHAN_RS[mst] ),  // 0 means no slice on channel - 1 means full slice on channel
            .ARCHAN_RS              ( MASTER_ARCHAN_RS[mst] ),  // 0 means no slice on channel - 1 means full slice on channel
            .RCHAN_RS               ( MASTER_RCHAN_RS[mst] ),    // 0 means no slice on channel - 1 means full slice on channel
            .WCHAN_RS               ( MASTER_WCHAN_RS[mst] ),    // 0 means no slice on channel - 1 means full slice on channel
            .BCHAN_RS               ( MASTER_BCHAN_RS[mst] ),    // 0 means no slice on channel - 1 means full slice on channel
            .OPEN_TRANS_MAX         ( OPEN_TRANS_MAX ),
            .ID_WIDTH               ( ID_WIDTH ), 
            .ADDR_WIDTH             ( ADDR_WIDTH ),
            .DATA_WIDTH             ( DATA_WIDTH ), 
            .MASTER_DATA_WIDTH      ( MASTER_PORTS_DATA_WIDTH[(mst+1)*32-1:mst*32] ),
	    .AHB_BRESP_CHECK_MODE          ( AHB_MASTER_PORTS_BRESP_CHECK_MODE[2*(mst+1)-1:2*mst] ),
	    .AHB_BRESP_CNT_WIDTH          ( AHB_MASTER_PORTS_BRESP_CNT_WIDTH[32*(mst+1)-1:32*mst] ),
            .SUPPORT_USER_SIGNALS   ( SUPPORT_USER_SIGNALS ),
            .USER_WIDTH             ( USER_WIDTH ),
            .CLOCK_DOMAIN_CROSSING  ( M_CDC[mst] )
          )
      mstrconv (
            // Global Signals
            .MST_CLK   ( M_CLK[mst] ),
            .XBAR_CLK  ( ACLK ),
            .ARESETN   ( ARESETN ),        // active low reset synchronoise to RE AClk - asserted async.
			.ACLK_syncReset (ACLK_syncReset),
    
            // Master Read Address Ports
            .MASTER_ARID       ( MASTER_ARID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH] ),
            .MASTER_ARADDR     ( MASTER_ARADDR[(mst+1)*ADDR_WIDTH-1:mst*ADDR_WIDTH] ),
            .MASTER_ARLEN      ( MASTER_ARLEN[(mst+1)*8-1:mst*8] ),
            .MASTER_ARSIZE     ( MASTER_ARSIZE[(mst+1)*3-1:mst*3] ),
            .MASTER_ARBURST    ( MASTER_ARBURST[(mst+1)*2-1:mst*2] ),
            .MASTER_ARLOCK     ( MASTER_ARLOCK[(mst+1)*2-1:mst*2] ),
            .MASTER_ARCACHE    ( MASTER_ARCACHE[(mst+1)*4-1:mst*4] ),
            .MASTER_ARPROT     ( MASTER_ARPROT[(mst+1)*3-1:mst*3]  ),
            .MASTER_ARREGION   ( MASTER_ARREGION[(mst+1)*4-1:mst*4] ),
            .MASTER_ARQOS      ( MASTER_ARQOS[(mst+1)*4-1:mst*4] ),
            .MASTER_ARUSER     ( MASTER_ARUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH] ),
            .MASTER_ARVALID    ( MASTER_ARVALID[mst] ),
            .MASTER_AWQOS      ( MASTER_AWQOS[(mst+1)*4-1:mst*4] ),
            .MASTER_AWREGION   ( MASTER_AWREGION[(mst+1)*4-1:mst*4] ),
            .MASTER_AWID       ( MASTER_AWID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH] ),
            .MASTER_AWADDR     ( MASTER_AWADDR[(mst+1)*ADDR_WIDTH-1:mst*ADDR_WIDTH] ),
            .MASTER_AWLEN      ( MASTER_AWLEN[(mst+1)*8-1:mst*8] ),
            .MASTER_AWSIZE     ( MASTER_AWSIZE[(mst+1)*3-1:mst*3] ),
            .MASTER_AWBURST    ( MASTER_AWBURST[(mst+1)*2-1:mst*2] ),
            .MASTER_AWLOCK     ( MASTER_AWLOCK[(mst+1)*2-1:mst*2] ),
            .MASTER_AWCACHE    ( MASTER_AWCACHE[(mst+1)*4-1:mst*4] ),
            .MASTER_AWPROT     ( MASTER_AWPROT[(mst+1)*3-1:mst*3] ),
            .MASTER_AWUSER     ( MASTER_AWUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH] ),
            .MASTER_AWVALID    ( MASTER_AWVALID[mst] ),
            .MASTER_WID        ( {ID_WIDTH{1'b0}} ),                           // jhayes : not used below currently, connected to avoid synthesis warning around unconnected mstnput.
            .MASTER_WDATA      ( MASTER_WDATA[MDW_UPPER_VEC[(1+mst)*13-1:13*mst]-1:MDW_LOWER_VEC[(1+mst)*13-1:13*mst]] ),
            .MASTER_WSTRB      ( MASTER_WSTRB[MDW_UPPER_VEC[(1+mst)*13-1:13*mst]/8-1:MDW_LOWER_VEC[(1+mst)*13-1:13*mst]/8] ),
            .MASTER_WLAST      ( MASTER_WLAST[mst] ),
            .MASTER_WUSER      ( MASTER_WUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH] ),
            .MASTER_WVALID     ( MASTER_WVALID[mst] ),
            .MASTER_BREADY     ( MASTER_BREADY[mst] ),
            .MASTER_RREADY     ( MASTER_RREADY[mst] ),
            .MASTER_ARREADY    ( MASTER_ARREADY[mst]),
            .MASTER_RID        ( MASTER_RID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH]),
            .MASTER_RDATA      ( MASTER_RDATA[MDW_UPPER_VEC[(1+mst)*13-1:13*mst]-1:MDW_LOWER_VEC[(1+mst)*13-1:13*mst]]),
            .MASTER_RRESP      ( MASTER_RRESP[(mst+1)*2-1:mst*2]),
            .MASTER_RUSER      ( MASTER_RUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH]),
            .MASTER_BID        ( MASTER_BID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH]),
            .MASTER_BRESP      ( MASTER_BRESP[(mst+1)*2-1:mst*2]),
            .MASTER_BUSER      ( MASTER_BUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH]),
            .MASTER_RLAST      ( MASTER_RLAST[mst]),
            .MASTER_RVALID     ( MASTER_RVALID[mst]),
            .MASTER_AWREADY    ( MASTER_AWREADY[mst]),
            .MASTER_WREADY     ( MASTER_WREADY[mst]),
            .MASTER_BVALID     ( MASTER_BVALID[mst]),

            .MASTER_HADDR          ( MASTER_HADDR[(mst+1)*32-1:mst*32] ),
            .MASTER_HBURST         ( MASTER_HBURST[(mst+1)*3-1:mst*3] ),
            .MASTER_HMASTLOCK      ( MASTER_HMASTLOCK[mst] ),
            .MASTER_HPROT          ( MASTER_HPROT[(mst+1)*7-1:mst*7] ),          
            .MASTER_HSIZE          ( MASTER_HSIZE[(mst+1)*3-1:mst*3] ),
            .MASTER_HNONSEC        ( MASTER_HNONSEC[mst] ),
            .MASTER_HTRANS         ( MASTER_HTRANS[(mst+1)*2-1:mst*2] ),
            .MASTER_HWDATA         ( MASTER_HWDATA[MDW_UPPER_VEC[(1+mst)*13-1:13*mst]-1:MDW_LOWER_VEC[(1+mst)*13-1:13*mst]] ),
            .MASTER_HRDATA         ( MASTER_HRDATA[MDW_UPPER_VEC[(1+mst)*13-1:13*mst]-1:MDW_LOWER_VEC[(1+mst)*13-1:13*mst]] ),
            .MASTER_HWRITE         ( MASTER_HWRITE[mst] ),
            .MASTER_HREADY         ( MASTER_HREADY[mst] ),
            .MASTER_HRESP          ( MASTER_HRESP[mst] ),
//            .MASTER_HEXOKAY      ( MASTER_HEXOKAY[mst] ),
//            .MASTER_HEXCL        ( MASTER_HEXCL[mst] ),
            .MASTER_HSEL           ( MASTER_HSEL[mst] ),

            .int_masterARID        ( masterARID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH] ),
            .int_masterARADDR      ( masterARADDR[(mst+1)*ADDR_WIDTH-1:mst*ADDR_WIDTH] ),
            .int_masterARLEN       ( masterARLEN[(mst+1)*8-1:mst*8] ),
            .int_masterARSIZE      ( masterARSIZE[(mst+1)*3-1:mst*3] ),
            .int_masterARBURST     ( masterARBURST[(mst+1)*2-1:mst*2] ),
            .int_masterARLOCK      ( masterARLOCK[(mst+1)*2-1:mst*2] ),
            .int_masterARCACHE     ( masterARCACHE[(mst+1)*4-1:mst*4] ),
            .int_masterARPROT      ( masterARPROT[(mst+1)*3-1:mst*3]  ),
            .int_masterARREGION    ( masterARREGION[(mst+1)*4-1:mst*4] ),
            .int_masterARQOS       ( masterARQOS[(mst+1)*4-1:mst*4] ),
            .int_masterARUSER      ( masterARUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH] ),
            .int_masterARVALID     ( masterARVALID[mst] ),
            .int_masterAWQOS       ( masterAWQOS[(mst+1)*4-1:mst*4] ),
            .int_masterAWREGION    ( masterAWREGION[(mst+1)*4-1:mst*4] ),
            .int_masterAWID        ( masterAWID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH] ),
            .int_masterAWADDR      ( masterAWADDR[(mst+1)*ADDR_WIDTH-1:mst*ADDR_WIDTH] ),
            .int_masterAWLEN       ( masterAWLEN[(mst+1)*8-1:mst*8] ),
            .int_masterAWSIZE      ( masterAWSIZE[(mst+1)*3-1:mst*3] ),
            .int_masterAWBURST     ( masterAWBURST[(mst+1)*2-1:mst*2] ),
            .int_masterAWLOCK      ( masterAWLOCK[(mst+1)*2-1:mst*2] ),
            .int_masterAWCACHE     ( masterAWCACHE[(mst+1)*4-1:mst*4] ),
            .int_masterAWPROT      ( masterAWPROT[(mst+1)*3-1:mst*3] ),
            .int_masterAWUSER      ( masterAWUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH] ),
            .int_masterAWVALID     ( masterAWVALID[mst] ),
            .int_masterWDATA       ( masterWDATA[(mst+1)*DATA_WIDTH-1:mst*DATA_WIDTH] ),
            .int_masterWSTRB       ( masterWSTRB[(mst+1)*DATA_WIDTH/8-1:mst*DATA_WIDTH/8] ),
            .int_masterWLAST       ( masterWLAST[mst] ),
            .int_masterWUSER       ( masterWUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH] ),
            .int_masterWVALID      ( masterWVALID[mst] ),
            .int_masterBREADY      ( masterBREADY[mst] ),
            .int_masterRREADY      ( masterRREADY[mst] ),
            .int_masterARREADY     ( masterARREADY[mst]),
            .int_masterRID         ( masterRID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH]),
            .int_masterRDATA       ( masterRDATA[(mst+1)*DATA_WIDTH-1:mst*DATA_WIDTH]),
            .int_masterRRESP       ( masterRRESP[(mst+1)*2-1:mst*2]),
            .int_masterRUSER       ( masterRUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH]),
            .int_masterBID         ( masterBID[(mst+1)*ID_WIDTH-1:mst*ID_WIDTH]),
            .int_masterBRESP       ( masterBRESP[(mst+1)*2-1:mst*2]),
            .int_masterBUSER       ( masterBUSER[(mst+1)*USER_WIDTH-1:mst*USER_WIDTH]),
            .int_masterRLAST       ( masterRLAST[mst]),
            .int_masterRVALID      ( masterRVALID[mst]),
            .int_masterAWREADY     ( masterAWREADY[mst]),
            .int_masterWREADY      ( masterWREADY[mst]),
            .int_masterBVALID      ( masterBVALID[mst])

          );
          end // MstConvertor_loop
  endgenerate   
  
   //===============================================================================================================================

        genvar slv;
  generate
                for (slv=0; slv<NUM_SLAVES; slv=slv+1) begin : SlvConvertor_loop
        caxi4interconnect_SlaveConvertor #
         (
              .SLAVE_TYPE            ( SLAVE_TYPE [(slv+1)*2-1:slv*2] ),  // Protocol type = AXI4 - 2'b00, AXI4Lite - 2'b01, AXI3 - 2'b10
              .DWC_DATA_FIFO_DEPTH   ( SLAVE_DWC_DATA_FIFO_DEPTH[(slv+1)*14-1:slv*14] ),
              .DWC_ADDR_FIFO_DEPTH_CEILING (DWC_ADDR_FIFO_DEPTH_CEILING),
              .SLAVE_NUMBER          ( slv ),          // master number
              .AWCHAN_RS             ( SLAVE_AWCHAN_RS[slv] ),  // 0 means no slice on channel - 1 means full slice on channel
              .ARCHAN_RS             ( SLAVE_ARCHAN_RS[slv] ),  // 0 means no slice on channel - 1 means full slice on channel
              .RCHAN_RS              ( SLAVE_RCHAN_RS[slv] ),  // 0 means no slice on channel - 1 means full slice on channel
              .WCHAN_RS              ( SLAVE_WCHAN_RS[slv] ),  // 0 means no slice on channel - 1 means full slice on channel
              .BCHAN_RS              ( SLAVE_BCHAN_RS[slv] ),  // 0 means no slice on channel - 1 means full slice on channel  
              .OPEN_TRANS_MAX        ( OPEN_TRANS_MAX ),
              .ID_WIDTH              ( NUM_MASTERS_WIDTH + ID_WIDTH ),    // includes infrastructure ID
              .ADDR_WIDTH            ( ADDR_WIDTH ),        
              .DATA_WIDTH            ( DATA_WIDTH ), 
              .SLAVE_DATA_WIDTH      (SLAVE_PORTS_DATA_WIDTH[(slv+1)*32-1:slv*32] ),
              .READ_ZERO_SLAVE_ID( SLAVE_READ_ZERO_SLAVE_ID[slv] & (SLAVE_PORTS_DATA_WIDTH[(slv+1)*32-1:slv*32] == DATA_WIDTH) ),
              .WRITE_ZERO_SLAVE_ID( SLAVE_WRITE_ZERO_SLAVE_ID[slv] & (SLAVE_PORTS_DATA_WIDTH[(slv+1)*32-1:slv*32] == DATA_WIDTH) ),
              .USER_WIDTH            ( USER_WIDTH ),
              .SLV_AXI4PRT_ADDRDEPTH ( SLV_AXI4PRT_ADDRDEPTH ),  // Number transations width - 1 => 2 transations, 2 => 4 transations, etc.
              .SLV_AXI4PRT_DATADEPTH ( SLV_AXI4PRT_DATADEPTH ),  // Number transations width - 1 => 2 transations, 2 => 4 transations, etc.
              .CLOCK_DOMAIN_CROSSING (S_CDC[slv])
          )
        slvcnv (
              .SLV_CLK  ( S_CLK[slv] ),
              .XBAR_CLK ( ACLK ),
              .ARESETN  ( ARESETN ),        // active low reset synchronoise to RE AClk - asserted async.
			  .ACLK_syncReset (ACLK_syncReset),
       
              .SLAVE_AWID        ( SLAVE_AWID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .SLAVE_AWADDR      ( SLAVE_AWADDR[(slv+1)*ADDR_WIDTH-1:slv*ADDR_WIDTH] ),  
              .SLAVE_AWLEN       ( SLAVE_AWLEN[(slv+1)*8-1:slv*8] ),  
              .SLAVE_AWSIZE      ( SLAVE_AWSIZE[(slv+1)*3-1:slv*3] ),  
              .SLAVE_AWBURST     ( SLAVE_AWBURST[(slv+1)*2-1:slv*2] ),  
              .SLAVE_AWLOCK      ( SLAVE_AWLOCK[(slv+1)*2-1:slv*2] ),  
              .SLAVE_AWCACHE     ( SLAVE_AWCACHE[(slv+1)*4-1:slv*4] ),  
              .SLAVE_AWPROT      ( SLAVE_AWPROT[(slv+1)*3-1:slv*3] ),  
              .SLAVE_AWREGION    ( SLAVE_AWREGION[(slv+1)*4-1:slv*4] ),   
              .SLAVE_AWQOS       ( SLAVE_AWQOS[(slv+1)*4-1:slv*4] ),  
              .SLAVE_AWUSER      ( SLAVE_AWUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .SLAVE_AWVALID     ( SLAVE_AWVALID[slv] ),
              .SLAVE_WID         ( SLAVE_WID[ (slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)]  ),
              .SLAVE_WDATA       ( SLAVE_WDATA[SDW_UPPER_VEC[(1+slv)*13-1:13*slv]-1:SDW_LOWER_VEC[(1+slv)*13-1:13*slv]] ),  
              .SLAVE_WSTRB       ( SLAVE_WSTRB[SDW_UPPER_VEC[(1+slv)*13-1:13*slv]/8-1:SDW_LOWER_VEC[(1+slv)*13-1:13*slv]/8] ),  
              .SLAVE_WLAST       ( SLAVE_WLAST[slv] ),  
              .SLAVE_WUSER       ( SLAVE_WUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .SLAVE_WVALID      ( SLAVE_WVALID[slv] ),      
              .SLAVE_BREADY      ( SLAVE_BREADY[slv] ),        
              .SLAVE_ARID        ( SLAVE_ARID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .SLAVE_ARADDR      ( SLAVE_ARADDR[(slv+1)*ADDR_WIDTH-1:slv*ADDR_WIDTH] ),  
              .SLAVE_ARLEN       ( SLAVE_ARLEN[(slv+1)*8-1:slv*8] ),  
              .SLAVE_ARSIZE      ( SLAVE_ARSIZE[(slv+1)*3-1:slv*3] ),  
              .SLAVE_ARBURST     ( SLAVE_ARBURST[(slv+1)*2-1:slv*2] ),  
              .SLAVE_ARLOCK      ( SLAVE_ARLOCK[(slv+1)*2-1:slv*2] ),  
              .SLAVE_ARCACHE     ( SLAVE_ARCACHE[(slv+1)*4-1:slv*4] ),  
              .SLAVE_ARPROT      ( SLAVE_ARPROT[(slv+1)*3-1:slv*3] ),  
              .SLAVE_ARREGION    ( SLAVE_ARREGION[(slv+1)*4-1:slv*4] ),   
              .SLAVE_ARQOS       ( SLAVE_ARQOS[(slv+1)*4-1:slv*4] ),  
              .SLAVE_ARUSER      ( SLAVE_ARUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .SLAVE_ARVALID     ( SLAVE_ARVALID[slv] ),      
              .SLAVE_RREADY      ( SLAVE_RREADY[slv] ),    
              .SLAVE_AWREADY     ( SLAVE_AWREADY[slv] ),          
              .SLAVE_WREADY      ( SLAVE_WREADY[slv] ),        
              .SLAVE_BID         ( SLAVE_BID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .SLAVE_BRESP       ( SLAVE_BRESP[(slv+1)*2-1:slv*2] ),  
              .SLAVE_BUSER       ( SLAVE_BUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .SLAVE_BVALID      ( SLAVE_BVALID[slv] ),        
              .SLAVE_ARREADY     ( SLAVE_ARREADY[slv] ),        
              .SLAVE_RID         ( SLAVE_RID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .SLAVE_RDATA       ( SLAVE_RDATA[SDW_UPPER_VEC[(1+slv)*13-1:13*slv]-1:SDW_LOWER_VEC[(1+slv)*13-1:13*slv]] ),  // Input to this file
              .SLAVE_RRESP       ( SLAVE_RRESP[(slv+1)*2-1:slv*2] ),  
              .SLAVE_RLAST       ( SLAVE_RLAST[slv] ),  
              .SLAVE_RUSER       ( SLAVE_RUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .SLAVE_RVALID      ( SLAVE_RVALID[slv] ),

              .slaveAWID        ( slaveAWID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .slaveAWADDR      ( slaveAWADDR[(slv+1)*ADDR_WIDTH-1:slv*ADDR_WIDTH] ),  
              .slaveAWLEN       ( slaveAWLEN[(slv+1)*8-1:slv*8] ),  
              .slaveAWSIZE      ( slaveAWSIZE[(slv+1)*3-1:slv*3] ),  
              .slaveAWBURST     ( slaveAWBURST[(slv+1)*2-1:slv*2] ),  
              .slaveAWLOCK      ( slaveAWLOCK[(slv+1)*2-1:slv*2] ),  
              .slaveAWCACHE     ( slaveAWCACHE[(slv+1)*4-1:slv*4] ),  
              .slaveAWPROT      ( slaveAWPROT[(slv+1)*3-1:slv*3] ),  
              .slaveAWREGION    ( slaveAWREGION[(slv+1)*4-1:slv*4] ),   
              .slaveAWQOS       ( slaveAWQOS[(slv+1)*4-1:slv*4] ),  
              .slaveAWUSER      ( slaveAWUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .slaveAWVALID     ( slaveAWVALID[slv] ),        
              .slaveWDATA       ( slaveWDATA[(slv+1)*DATA_WIDTH-1:slv*DATA_WIDTH] ),  
              .slaveWSTRB       ( slaveWSTRB[(slv+1)*DATA_WIDTH/8-1:slv*DATA_WIDTH/8] ),  
              .slaveWLAST       ( slaveWLAST[slv] ),  
              .slaveWUSER       ( slaveWUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .slaveWVALID      ( slaveWVALID[slv] ),      
              .slaveBREADY      ( slaveBREADY[slv] ),        
              .slaveARID        ( slaveARID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .slaveARADDR      ( slaveARADDR[(slv+1)*ADDR_WIDTH-1:slv*ADDR_WIDTH] ),  
              .slaveARLEN       ( slaveARLEN[(slv+1)*8-1:slv*8] ),  
              .slaveARSIZE      ( slaveARSIZE[(slv+1)*3-1:slv*3] ),  
              .slaveARBURST     ( slaveARBURST[(slv+1)*2-1:slv*2] ),  
              .slaveARLOCK      ( slaveARLOCK[(slv+1)*2-1:slv*2] ),  
              .slaveARCACHE     ( slaveARCACHE[(slv+1)*4-1:slv*4] ),  
              .slaveARPROT      ( slaveARPROT[(slv+1)*3-1:slv*3] ),  
              .slaveARREGION    ( slaveARREGION[(slv+1)*4-1:slv*4] ),   
              .slaveARQOS       ( slaveARQOS[(slv+1)*4-1:slv*4] ),  
              .slaveARUSER      ( slaveARUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .slaveARVALID     ( slaveARVALID[slv] ),      
              .slaveRREADY      ( slaveRREADY[slv] ),        
              .slaveAWREADY     ( slaveAWREADY[slv] ),          
              .slaveWREADY      ( slaveWREADY[slv] ),        
              .slaveBID         ( slaveBID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .slaveBRESP       ( slaveBRESP[(slv+1)*2-1:slv*2] ),  
              .slaveBUSER       ( slaveBUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .slaveBVALID      ( slaveBVALID[slv] ),        
              .slaveARREADY     ( slaveARREADY[slv] ),        
              .slaveRID         ( slaveRID[(slv+1)*(NUM_MASTERS_WIDTH+ID_WIDTH)-1:slv*(NUM_MASTERS_WIDTH+ID_WIDTH)] ),  
              .slaveRDATA       ( slaveRDATA[(slv+1)*DATA_WIDTH-1:slv*DATA_WIDTH] ),  // Output from this module, input to this file
              .slaveRRESP       ( slaveRRESP[(slv+1)*2-1:slv*2] ),  
              .slaveRLAST       ( slaveRLAST[slv] ),  
              .slaveRUSER       ( slaveRUSER[(slv+1)*USER_WIDTH-1:slv*USER_WIDTH] ),  
              .slaveRVALID      ( slaveRVALID[slv] )
            ); 
    end //SlvConvertor_loop
  endgenerate     
endmodule  // COREAXI4INTERCONNECT.v
