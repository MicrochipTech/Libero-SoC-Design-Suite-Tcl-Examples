// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAOI00
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAOO1
,
CAXI4DMAIO1
,
CAXI4DMAIlOl
,
CAXI4DMAlO1
,
CAXI4DMAIO1l
,
CAXI4DMAlI1
,
CAXI4DMAII00
,
CAXI4DMAlI00
,
CAXI4DMAOl00
,
CAXI4DMAlOO0
,
CAXI4DMAI1Il
,
CAXI4DMAIl00
,
CAXI4DMAll00
)
;
parameter
CAXI4DMAO000
=
1
;
parameter
CAXI4DMAI000
=
1
;
function
integer
CAXI4DMAIOII
;
input
integer
CAXI4DMAlOII
;
integer
CAXI4DMAOIII
,
CAXI4DMAIIII
,
CAXI4DMAlIII
;
begin
CAXI4DMAIIII
=
1
;
CAXI4DMAlIII
=
0
;
CAXI4DMAOIII
=
CAXI4DMAlOII
+
1
;
while
(
CAXI4DMAIIII
<
CAXI4DMAOIII
)
begin
CAXI4DMAIIII
=
CAXI4DMAIIII
*
2
;
CAXI4DMAlIII
=
CAXI4DMAlIII
+
1
;
end
CAXI4DMAIOII
=
CAXI4DMAlIII
;
end
endfunction
localparam
CAXI4DMAl000
=
CAXI4DMAI000
*
CAXI4DMAO000
;
localparam
CAXI4DMAOlII
=
CAXI4DMAIOII
(
CAXI4DMAO000
)
;
localparam
CAXI4DMAO100
=
CAXI4DMAIOII
(
CAXI4DMAl000
)
;
localparam
CAXI4DMAI100
=
CAXI4DMAIOII
(
CAXI4DMAI000
-
1
)
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAOO1
;
input
[
CAXI4DMAI100
-
1
:
0
]
CAXI4DMAIO1
;
input
[
(
CAXI4DMAO000
*
8
)
-
1
:
0
]
CAXI4DMAlO1
;
input
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAIlOl
;
input
CAXI4DMAIO1l
;
input
[
CAXI4DMAI100
-
1
:
0
]
CAXI4DMAlI1
;
input
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAII00
;
input
CAXI4DMAlI00
;
input
CAXI4DMAOl00
;
input
CAXI4DMAlOO0
;
output
[
(
CAXI4DMAO000
*
8
)
-
1
:
0
]
CAXI4DMAI1Il
;
output
[
CAXI4DMAO100
-
1
:
0
]
CAXI4DMAIl00
;
output
[
CAXI4DMAO100
-
1
:
0
]
CAXI4DMAll00
;
reg
[
(
CAXI4DMAO000
*
8
)
-
1
:
0
]
CAXI4DMAl100
[
0
:
CAXI4DMAI000
-
1
]
;
reg
[
(
CAXI4DMAO000
*
8
)
-
1
:
0
]
CAXI4DMAOO10
[
0
:
CAXI4DMAI000
-
1
]
;
reg
[
CAXI4DMAO100
-
1
:
0
]
CAXI4DMAIO10
;
reg
[
CAXI4DMAO100
-
1
:
0
]
CAXI4DMAlO10
;
wire
[
3
:
0
]
CAXI4DMAOI10
;
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAOO1
)
begin
if
(
CAXI4DMAOl00
)
begin
CAXI4DMAOO10
[
CAXI4DMAIO1
]
<=
CAXI4DMAlO1
;
end
else
begin
CAXI4DMAl100
[
CAXI4DMAIO1
]
<=
CAXI4DMAlO1
;
end
end
end
assign
CAXI4DMAI1Il
=
(
CAXI4DMAlI00
)
?
CAXI4DMAOO10
[
CAXI4DMAlI1
]
:
CAXI4DMAl100
[
CAXI4DMAlI1
]
;
assign
CAXI4DMAOI10
=
{
CAXI4DMAOO1
,
CAXI4DMAOl00
,
CAXI4DMAIO1l
,
CAXI4DMAlI00
}
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO10
<=
{
CAXI4DMAO100
{
1
'b
0
}
}
;
CAXI4DMAlO10
<=
{
CAXI4DMAO100
{
1
'b
0
}
}
;
end
else
begin
if
(
CAXI4DMAlOO0
)
begin
if
(
CAXI4DMAlI00
)
begin
CAXI4DMAlO10
<=
{
CAXI4DMAO100
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIO10
<=
{
CAXI4DMAO100
{
1
'b
0
}
}
;
end
if
(
(
CAXI4DMAOO1
==
1
'b
1
)
&&
(
CAXI4DMAlI00
!=
CAXI4DMAOl00
)
)
begin
if
(
CAXI4DMAOl00
)
begin
CAXI4DMAlO10
<=
CAXI4DMAlO10
+
CAXI4DMAIlOl
;
end
else
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
+
CAXI4DMAIlOl
;
end
end
end
else
begin
case
(
CAXI4DMAOI10
)
4
'b
0010
,
4
'b
0110
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
-
CAXI4DMAII00
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
;
end
4
'b
0011
,
4
'b
0111
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
-
CAXI4DMAII00
;
end
4
'b
1000
,
4
'b
1001
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
+
CAXI4DMAIlOl
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
;
end
4
'b
1010
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
+
CAXI4DMAIlOl
-
CAXI4DMAII00
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
;
end
4
'b
1011
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
+
CAXI4DMAIlOl
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
-
CAXI4DMAII00
;
end
4
'b
1100
,
4
'b
1101
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
+
CAXI4DMAIlOl
;
end
4
'b
1110
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
-
CAXI4DMAII00
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
+
CAXI4DMAIlOl
;
end
4
'b
1111
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
+
CAXI4DMAIlOl
-
CAXI4DMAII00
;
end
default
:
begin
CAXI4DMAIO10
<=
CAXI4DMAIO10
;
CAXI4DMAlO10
<=
CAXI4DMAlO10
;
end
endcase
end
end
end
assign
CAXI4DMAIl00
=
(
CAXI4DMAlI00
)
?
CAXI4DMAlO10
:
CAXI4DMAIO10
;
assign
CAXI4DMAll00
=
(
CAXI4DMAOl00
)
?
CAXI4DMAlO10
:
CAXI4DMAIO10
;
endmodule
