// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAOlIll
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAll1l
,
CAXI4DMAO01l
,
CAXI4DMAI01l
,
CAXI4DMAl01l
,
CAXI4DMAO11l
,
valid
,
CAXI4DMAlIlOI
,
CAXI4DMAOllOI
,
CAXI4DMAIllOI
,
CAXI4DMAOI0OI
,
intDscrptrNum
,
CAXI4DMAII0OI
,
CAXI4DMAlI0OI
,
strDscrptr
,
CAXI4DMAOIO0
,
CAXI4DMAO0Ill
,
CAXI4DMAI0Ill
)
;
parameter
CAXI4DMAIlIll
=
1
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAll1l
;
input
CAXI4DMAO01l
;
input
[
1
:
0
]
CAXI4DMAI01l
;
input
[
31
:
0
]
CAXI4DMAl01l
;
input
CAXI4DMAO11l
;
input
valid
;
input
CAXI4DMAlIlOI
;
input
CAXI4DMAOllOI
;
input
CAXI4DMAIllOI
;
input
CAXI4DMAOI0OI
;
input
[
4
:
0
]
intDscrptrNum
;
input
CAXI4DMAII0OI
;
input
[
31
:
0
]
CAXI4DMAlI0OI
;
input
strDscrptr
;
output
[
31
:
0
]
CAXI4DMAOIO0
;
output
CAXI4DMAO0Ill
;
output
reg
CAXI4DMAI0Ill
;
localparam
CAXI4DMAl0O0l
=
1
'b
0
;
localparam
CAXI4DMAO1O0l
=
1
'b
1
;
reg
CAXI4DMAl10OI
;
reg
CAXI4DMAOO1OI
;
wire
[
5
:
0
]
CAXI4DMAOIIll
;
wire
[
41
:
0
]
CAXI4DMAI1O0l
;
wire
[
41
:
0
]
CAXI4DMAl1O0l
;
wire
[
41
:
0
]
CAXI4DMAOOI0l
;
reg
CAXI4DMAIOI0l
;
wire
CAXI4DMAlOI0l
;
wire
CAXI4DMAO0Ill
;
wire
CAXI4DMAOII0l
;
wire
CAXI4DMAIII0l
;
wire
CAXI4DMAlII0l
;
wire
[
3
:
0
]
CAXI4DMAOlI0l
;
reg
[
3
:
0
]
CAXI4DMAIlI0l
;
reg
[
3
:
0
]
CAXI4DMAllI0l
;
reg
[
41
:
0
]
CAXI4DMAO0I0l
;
assign
CAXI4DMAOIIll
=
(
strDscrptr
)
?
6
'd
33
:
(
CAXI4DMAII0OI
)
?
6
'd
32
:
intDscrptrNum
;
assign
CAXI4DMAI1O0l
=
{
CAXI4DMAlI0OI
,
CAXI4DMAOIIll
,
CAXI4DMAOI0OI
,
CAXI4DMAIllOI
,
CAXI4DMAOllOI
,
CAXI4DMAlIlOI
}
;
CAXI4DMAII10
#
(
.CAXI4DMAll10
(
42
)
,
.CAXI4DMAO010
(
CAXI4DMAIlIll
)
)
CAXI4DMAI0I0l
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAOO1
(
valid
)
,
.CAXI4DMAlO1
(
CAXI4DMAI1O0l
)
,
.CAXI4DMAIO1l
(
CAXI4DMAlOI0l
)
,
.CAXI4DMAI1Il
(
CAXI4DMAOOI0l
)
,
.CAXI4DMAlI10
(
)
,
.CAXI4DMAOl10
(
CAXI4DMAO0Ill
)
,
.CAXI4DMAIl10
(
CAXI4DMAOII0l
)
)
;
assign
CAXI4DMAIII0l
=
!
CAXI4DMAOII0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAl0O0l
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
case
(
CAXI4DMAl10OI
)
CAXI4DMAl0O0l
:
begin
if
(
CAXI4DMAIII0l
)
begin
CAXI4DMAIOI0l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1O0l
;
end
else
begin
CAXI4DMAIOI0l
<=
1
'b
0
;
CAXI4DMAOO1OI
<=
CAXI4DMAl0O0l
;
end
end
CAXI4DMAO1O0l
:
begin
CAXI4DMAIOI0l
<=
1
'b
0
;
if
(
CAXI4DMAlOI0l
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl0O0l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1O0l
;
end
end
endcase
end
assign
CAXI4DMAlOI0l
=
~
CAXI4DMAlII0l
&
CAXI4DMAI0Ill
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAllI0l
<=
4
'b
0
;
end
else
begin
if
(
CAXI4DMAll1l
&
CAXI4DMAO01l
&
CAXI4DMAO11l
&&
(
CAXI4DMAI01l
[
1
:
0
]
==
2
'b
10
)
)
begin
CAXI4DMAllI0l
<=
CAXI4DMAl01l
[
3
:
0
]
;
end
else
begin
CAXI4DMAllI0l
<=
4
'b
0
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIlI0l
<=
4
'b
0
;
end
else
begin
if
(
CAXI4DMAll1l
&
CAXI4DMAO01l
&
CAXI4DMAO11l
&&
(
CAXI4DMAI01l
[
1
:
0
]
==
2
'b
01
)
)
begin
CAXI4DMAIlI0l
<=
CAXI4DMAl01l
[
3
:
0
]
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO0I0l
<=
42
'b
0
;
end
else
begin
if
(
CAXI4DMAIOI0l
)
begin
CAXI4DMAO0I0l
<=
CAXI4DMAOOI0l
[
41
:
0
]
;
end
else
begin
CAXI4DMAO0I0l
<=
{
CAXI4DMAO0I0l
[
41
:
4
]
,
CAXI4DMAl1O0l
[
3
:
0
]
}
;
end
end
end
assign
CAXI4DMAl1O0l
=
CAXI4DMAO0I0l
[
3
:
0
]
&
~
CAXI4DMAllI0l
[
3
:
0
]
;
assign
CAXI4DMAOlI0l
=
CAXI4DMAl1O0l
[
3
:
0
]
&
CAXI4DMAIlI0l
[
3
:
0
]
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI0Ill
<=
1
'b
0
;
end
else
begin
CAXI4DMAI0Ill
<=
CAXI4DMAlII0l
;
end
end
assign
CAXI4DMAlII0l
=
(
|
CAXI4DMAOlI0l
[
3
:
0
]
)
;
assign
CAXI4DMAOIO0
=
(
CAXI4DMAI01l
==
2
'b
11
)
?
CAXI4DMAO0I0l
[
41
:
10
]
:
(
CAXI4DMAI01l
==
2
'b
01
)
?
{
{
28
{
1
'b
0
}
}
,
CAXI4DMAIlI0l
[
3
:
0
]
}
:
(
CAXI4DMAI01l
==
2
'b
10
)
?
32
'b
0
:
{
{
22
{
1
'b
0
}
}
,
CAXI4DMAO0I0l
[
9
:
0
]
}
;
endmodule
