// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAI1OOI
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAll1
,
CAXI4DMAO01
,
CAXI4DMAl01
,
CAXI4DMAO11
,
CAXI4DMAI11
,
CAXI4DMAl11
,
CAXI4DMAIIOI
,
CAXI4DMAlIOI
,
CAXI4DMAOlOI
,
CAXI4DMAOOIOI
,
CAXI4DMAOIO0
,
CAXI4DMAIIO0
,
CAXI4DMAlOl
,
CAXI4DMAIIl
,
CAXI4DMAOll
,
CAXI4DMAIll
,
CAXI4DMAlll
,
CAXI4DMAO0l
,
CAXI4DMAI0l
,
CAXI4DMAl0l
,
CAXI4DMAll1l
,
CAXI4DMAO01l
,
CAXI4DMAI01l
,
CAXI4DMAl01l
,
CAXI4DMAO11l
)
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAll1
;
input
CAXI4DMAO01
;
input
CAXI4DMAl01
;
input
CAXI4DMAO11
;
input
CAXI4DMAI11
;
input
[
10
:
0
]
CAXI4DMAl11
;
input
[
3
:
0
]
CAXI4DMAIIOI
;
input
[
31
:
0
]
CAXI4DMAlIOI
;
input
[
10
:
0
]
CAXI4DMAOlOI
;
input
CAXI4DMAOOIOI
;
input
[
31
:
0
]
CAXI4DMAOIO0
;
input
CAXI4DMAIIO0
;
output
[
1
:
0
]
CAXI4DMAlOl
;
output
[
31
:
0
]
CAXI4DMAIIl
;
output
CAXI4DMAOll
;
output
CAXI4DMAIll
;
output
CAXI4DMAlll
;
output
CAXI4DMAO0l
;
output
CAXI4DMAI0l
;
output
[
1
:
0
]
CAXI4DMAl0l
;
output
CAXI4DMAll1l
;
output
CAXI4DMAO01l
;
output
[
10
:
0
]
CAXI4DMAI01l
;
output
[
31
:
0
]
CAXI4DMAl01l
;
output
[
3
:
0
]
CAXI4DMAO11l
;
reg
[
8
:
0
]
CAXI4DMAl10OI
;
reg
[
8
:
0
]
CAXI4DMAOO1OI
;
reg
[
1
:
0
]
CAXI4DMAIO1OI
;
reg
[
1
:
0
]
CAXI4DMAlO1OI
;
reg
[
31
:
0
]
CAXI4DMAOI1OI
;
reg
[
31
:
0
]
CAXI4DMAII1OI
;
reg
CAXI4DMAlI1OI
;
reg
CAXI4DMAOl1OI
;
reg
CAXI4DMAIl1OI
;
reg
CAXI4DMAll1OI
;
reg
CAXI4DMAO01OI
;
reg
CAXI4DMAI01OI
;
reg
CAXI4DMAl01OI
;
reg
CAXI4DMAO11OI
;
reg
CAXI4DMAI11OI
;
reg
CAXI4DMAl11OI
;
reg
[
1
:
0
]
CAXI4DMAOOOII
;
reg
[
1
:
0
]
CAXI4DMAIOOII
;
reg
CAXI4DMAlOOII
;
reg
CAXI4DMAOIOII
;
reg
CAXI4DMAIIOII
;
reg
CAXI4DMAlIOII
;
reg
[
10
:
0
]
CAXI4DMAOlOII
;
reg
[
10
:
0
]
CAXI4DMAIlOII
;
reg
[
31
:
0
]
CAXI4DMAllOII
;
reg
[
31
:
0
]
CAXI4DMAO0OII
;
reg
[
3
:
0
]
CAXI4DMAI0OII
;
reg
[
3
:
0
]
CAXI4DMAl0OII
;
localparam
[
8
:
0
]
CAXI4DMAO1OII
=
9
'b
000000001
;
localparam
[
8
:
0
]
CAXI4DMAI1OII
=
9
'b
000000010
;
localparam
[
8
:
0
]
CAXI4DMAl1OII
=
9
'b
000000100
;
localparam
[
8
:
0
]
CAXI4DMAOOIII
=
9
'b
000001000
;
localparam
[
8
:
0
]
CAXI4DMAIOIII
=
9
'b
000010000
;
localparam
[
8
:
0
]
CAXI4DMAlOIII
=
9
'b
000100000
;
localparam
[
8
:
0
]
CAXI4DMAOIIII
=
9
'b
001000000
;
localparam
[
8
:
0
]
CAXI4DMAIIIII
=
9
'b
010000000
;
localparam
[
8
:
0
]
CAXI4DMAlIIII
=
9
'b
100000000
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAOl1OI
<=
1
'b
0
;
CAXI4DMAlO1OI
<=
2
'b
0
;
CAXI4DMAII1OI
<=
CAXI4DMAOI1OI
;
CAXI4DMAOl1OI
<=
1
'b
0
;
CAXI4DMAll1OI
<=
1
'b
0
;
CAXI4DMAI01OI
<=
1
'b
0
;
CAXI4DMAO11OI
<=
1
'b
0
;
CAXI4DMAl11OI
<=
1
'b
0
;
CAXI4DMAIOOII
<=
2
'b
0
;
CAXI4DMAOIOII
<=
CAXI4DMAlOOII
;
CAXI4DMAlIOII
<=
CAXI4DMAIIOII
;
CAXI4DMAIlOII
<=
CAXI4DMAOlOII
;
CAXI4DMAO0OII
<=
CAXI4DMAllOII
;
CAXI4DMAl0OII
<=
CAXI4DMAI0OII
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAll1
)
begin
CAXI4DMAOl1OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI1OII
;
end
else
if
(
CAXI4DMAO11
)
begin
CAXI4DMAO11OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOIIII
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAI1OII
:
begin
if
(
CAXI4DMAll1
&
CAXI4DMAOll
)
begin
CAXI4DMAIlOII
<=
{
CAXI4DMAl11
[
10
:
2
]
,
{
2
{
1
'b
0
}
}
}
;
if
(
CAXI4DMAO01
)
begin
CAXI4DMAOIOII
<=
1
'b
1
;
CAXI4DMAlIOII
<=
1
'b
1
;
CAXI4DMAO0OII
<=
CAXI4DMAlIOI
;
CAXI4DMAl0OII
<=
CAXI4DMAIIOI
;
CAXI4DMAOO1OI
<=
CAXI4DMAOOIII
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl1OII
;
end
end
else
begin
CAXI4DMAOl1OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI1OII
;
end
end
CAXI4DMAl1OII
:
begin
if
(
CAXI4DMAO01
)
begin
CAXI4DMAOIOII
<=
1
'b
1
;
CAXI4DMAlIOII
<=
1
'b
1
;
CAXI4DMAO0OII
<=
CAXI4DMAlIOI
;
CAXI4DMAl0OII
<=
CAXI4DMAIIOI
;
CAXI4DMAOO1OI
<=
CAXI4DMAOOIII
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl1OII
;
end
end
CAXI4DMAOOIII
:
begin
if
(
CAXI4DMAOOIOI
)
begin
CAXI4DMAIlOII
<=
11
'b
0
;
CAXI4DMAOIOII
<=
1
'b
0
;
CAXI4DMAlIOII
<=
1
'b
0
;
CAXI4DMAO0OII
<=
32
'b
0
;
CAXI4DMAl0OII
<=
4
'b
0
;
CAXI4DMAll1OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIOIII
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOOIII
;
end
end
CAXI4DMAIOIII
:
begin
if
(
CAXI4DMAIll
&
CAXI4DMAO01
)
begin
CAXI4DMAI01OI
<=
1
'b
1
;
CAXI4DMAlO1OI
<=
2
'b
00
;
CAXI4DMAOO1OI
<=
CAXI4DMAlOIII
;
end
else
begin
CAXI4DMAll1OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIOIII
;
end
end
CAXI4DMAlOIII
:
begin
if
(
CAXI4DMAl01
&
CAXI4DMAlll
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAI01OI
<=
1
'b
1
;
CAXI4DMAlO1OI
<=
2
'b
00
;
CAXI4DMAOO1OI
<=
CAXI4DMAlOIII
;
end
end
CAXI4DMAOIIII
:
begin
if
(
CAXI4DMAO11
&
CAXI4DMAO0l
)
begin
CAXI4DMAIlOII
<=
{
CAXI4DMAOlOI
[
10
:
2
]
,
{
2
{
1
'b
0
}
}
}
;
CAXI4DMAOIOII
<=
1
'b
1
;
CAXI4DMAlIOII
<=
1
'b
0
;
CAXI4DMAOO1OI
<=
CAXI4DMAIIIII
;
end
else
begin
CAXI4DMAO11OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOIIII
;
end
end
CAXI4DMAIIIII
:
begin
if
(
CAXI4DMAIIO0
)
begin
CAXI4DMAIlOII
<=
11
'b
0
;
CAXI4DMAIOOII
<=
2
'b
00
;
CAXI4DMAl11OI
<=
1
'b
1
;
CAXI4DMAII1OI
<=
CAXI4DMAOIO0
;
CAXI4DMAOO1OI
<=
CAXI4DMAlIIII
;
end
else
begin
CAXI4DMAOIOII
<=
1
'b
1
;
CAXI4DMAlIOII
<=
1
'b
0
;
CAXI4DMAOO1OI
<=
CAXI4DMAIIIII
;
end
end
CAXI4DMAlIIII
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
)
begin
CAXI4DMAII1OI
<=
32
'b
0
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAIOOII
<=
2
'b
00
;
CAXI4DMAl11OI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlIIII
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI1OI
<=
1
'b
0
;
end
else
begin
CAXI4DMAlI1OI
<=
CAXI4DMAOl1OI
;
end
end
assign
CAXI4DMAOll
=
CAXI4DMAlI1OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl01OI
<=
1
'b
0
;
end
else
begin
CAXI4DMAl01OI
<=
CAXI4DMAO11OI
;
end
end
assign
CAXI4DMAO0l
=
CAXI4DMAl01OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOI1OI
<=
32
'b
0
;
end
else
begin
CAXI4DMAOI1OI
<=
CAXI4DMAII1OI
;
end
end
assign
CAXI4DMAIIl
=
CAXI4DMAOI1OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIl1OI
<=
1
'b
0
;
end
else
begin
CAXI4DMAIl1OI
<=
CAXI4DMAll1OI
;
end
end
assign
CAXI4DMAIll
=
CAXI4DMAIl1OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO01OI
<=
1
'b
0
;
end
else
begin
CAXI4DMAO01OI
<=
CAXI4DMAI01OI
;
end
end
assign
CAXI4DMAlll
=
CAXI4DMAO01OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO1OI
<=
2
'b
0
;
end
else
begin
CAXI4DMAIO1OI
<=
CAXI4DMAlO1OI
;
end
end
assign
CAXI4DMAlOl
=
CAXI4DMAIO1OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI11OI
<=
1
'b
0
;
end
else
begin
CAXI4DMAI11OI
<=
CAXI4DMAl11OI
;
end
end
assign
CAXI4DMAI0l
=
CAXI4DMAI11OI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOOOII
<=
2
'b
0
;
end
else
begin
CAXI4DMAOOOII
<=
CAXI4DMAIOOII
;
end
end
assign
CAXI4DMAl0l
=
CAXI4DMAOOOII
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlOOII
<=
1
'b
0
;
end
else
begin
CAXI4DMAlOOII
<=
CAXI4DMAOIOII
;
end
end
assign
CAXI4DMAll1l
=
CAXI4DMAlOOII
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIIOII
<=
1
'b
0
;
end
else
begin
CAXI4DMAIIOII
<=
CAXI4DMAlIOII
;
end
end
assign
CAXI4DMAO01l
=
CAXI4DMAIIOII
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOlOII
<=
11
'b
0
;
end
else
begin
CAXI4DMAOlOII
<=
CAXI4DMAIlOII
;
end
end
assign
CAXI4DMAI01l
=
CAXI4DMAOlOII
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAllOII
<=
32
'b
0
;
end
else
begin
CAXI4DMAllOII
<=
CAXI4DMAO0OII
;
end
end
assign
CAXI4DMAl01l
=
CAXI4DMAllOII
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI0OII
<=
4
'b
0
;
end
else
begin
CAXI4DMAI0OII
<=
CAXI4DMAl0OII
;
end
end
assign
CAXI4DMAO11l
=
CAXI4DMAI0OII
;
endmodule
