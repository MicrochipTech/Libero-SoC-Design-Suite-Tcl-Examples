// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAIOI0I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAl0IlI
,
CAXI4DMAO1IlI
,
CAXI4DMAOII0I
,
CAXI4DMAIII0I
,
CAXI4DMAlII0I
,
CAXI4DMAOI0lI
,
CAXI4DMAOIllI
,
CAXI4DMAl1IlI
,
CAXI4DMAOOllI
,
CAXI4DMAIOllI
,
CAXI4DMAlI0OI
,
CAXI4DMAO1IOI
,
CAXI4DMAOlI0I
,
CAXI4DMAIIllI
,
CAXI4DMAIlI0I
,
CAXI4DMAlI0lI
,
CAXI4DMAlll1
)
;
parameter
CAXI4DMAlI1lI
=
4
;
parameter
CAXI4DMAOl1lI
=
2
;
parameter
CAXI4DMAl0OI
=
24
;
parameter
CAXI4DMAl1OI
=
133
;
parameter
CAXI4DMAO1llI
=
(
CAXI4DMAl1OI
+
1
+
32
)
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAl0IlI
;
input
CAXI4DMAO1IlI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAOII0I
;
input
CAXI4DMAIII0I
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAlII0I
;
input
CAXI4DMAOI0lI
;
input
CAXI4DMAOIllI
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl1IlI
;
input
[
31
:
0
]
CAXI4DMAOOllI
;
input
[
31
:
0
]
CAXI4DMAIOllI
;
input
[
31
:
0
]
CAXI4DMAlI0OI
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAOlI0I
;
input
CAXI4DMAIIllI
;
output
[
CAXI4DMAO1llI
-
1
:
0
]
CAXI4DMAIlI0I
;
output
reg
[
CAXI4DMAlI1lI
-
1
:
0
]
CAXI4DMAlI0lI
;
output
reg
[
CAXI4DMAlI1lI
-
1
:
0
]
CAXI4DMAlll1
;
reg
[
12
:
0
]
CAXI4DMAIIO0l
[
0
:
CAXI4DMAlI1lI
-
1
]
;
reg
[
63
:
0
]
CAXI4DMAlIO0l
[
0
:
CAXI4DMAlI1lI
-
1
]
;
reg
[
87
:
0
]
CAXI4DMAOlO0l
[
0
:
CAXI4DMAlI1lI
-
1
]
;
reg
[
CAXI4DMAlI1lI
-
1
:
0
]
CAXI4DMAIlO0l
;
integer
CAXI4DMAllO0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
CAXI4DMAlI0lI
<=
{
CAXI4DMAlI1lI
{
1
'b
0
}
}
;
else
if
(
CAXI4DMAl0IlI
&
!
CAXI4DMAO1IlI
)
CAXI4DMAlI0lI
[
CAXI4DMAOII0I
]
<=
CAXI4DMAIII0I
;
else
if
(
CAXI4DMAOI0lI
&&
!
CAXI4DMAOIllI
&&
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
)
CAXI4DMAlI0lI
[
CAXI4DMAlII0I
]
<=
1
'b
0
;
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
CAXI4DMAIlO0l
<=
{
CAXI4DMAlI1lI
{
1
'b
0
}
}
;
else
if
(
CAXI4DMAl0IlI
&
!
CAXI4DMAO1IlI
&
CAXI4DMAIII0I
)
CAXI4DMAIlO0l
[
CAXI4DMAOII0I
]
<=
CAXI4DMAO1IOI
[
13
]
;
else
if
(
CAXI4DMAOI0lI
&&
!
CAXI4DMAOIllI
&&
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
)
CAXI4DMAIlO0l
[
CAXI4DMAlII0I
]
<=
1
'b
0
;
else
if
(
CAXI4DMAOI0lI
&
!
CAXI4DMAOIllI
&
CAXI4DMAIIllI
)
CAXI4DMAIlO0l
[
CAXI4DMAlII0I
]
<=
1
'b
1
;
end
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAl0IlI
&
!
CAXI4DMAO1IlI
)
CAXI4DMAlIO0l
[
CAXI4DMAOII0I
]
<=
{
CAXI4DMAlI0OI
,
CAXI4DMAO1IOI
[
133
:
102
]
}
;
end
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAl0IlI
&
!
CAXI4DMAO1IlI
)
CAXI4DMAIIO0l
[
CAXI4DMAOII0I
]
<=
CAXI4DMAO1IOI
[
12
:
0
]
;
end
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAl0IlI
&
!
CAXI4DMAO1IlI
)
CAXI4DMAOlO0l
[
CAXI4DMAOII0I
]
<=
CAXI4DMAO1IOI
[
101
:
14
]
;
else
if
(
CAXI4DMAOI0lI
&
!
CAXI4DMAOIllI
)
CAXI4DMAOlO0l
[
CAXI4DMAlII0I
]
<=
{
CAXI4DMAIOllI
,
CAXI4DMAOOllI
,
CAXI4DMAl1IlI
}
;
end
assign
CAXI4DMAIlI0I
=
{
CAXI4DMAlI0lI
[
CAXI4DMAOlI0I
]
,
CAXI4DMAlIO0l
[
CAXI4DMAOlI0I
]
,
CAXI4DMAOlO0l
[
CAXI4DMAOlI0I
]
,
CAXI4DMAIlO0l
[
CAXI4DMAOlI0I
]
,
CAXI4DMAIIO0l
[
CAXI4DMAOlI0I
]
}
;
always
@
(
*
)
begin
for
(
CAXI4DMAllO0l
=
0
;
CAXI4DMAllO0l
<=
CAXI4DMAlI1lI
-
1
;
CAXI4DMAllO0l
=
CAXI4DMAllO0l
+
1
)
begin
if
(
(
CAXI4DMAllO0l
==
CAXI4DMAlII0I
)
&&
!
CAXI4DMAlI0lI
[
CAXI4DMAllO0l
]
)
begin
CAXI4DMAlll1
[
CAXI4DMAllO0l
]
=
(
CAXI4DMAOI0lI
&&
!
CAXI4DMAOIllI
&&
(
CAXI4DMAl1IlI
==
{
CAXI4DMAl0OI
{
1
'b
0
}
}
)
)
;
end
else
begin
CAXI4DMAlll1
[
CAXI4DMAllO0l
]
=
1
'b
0
;
end
end
end
endmodule
