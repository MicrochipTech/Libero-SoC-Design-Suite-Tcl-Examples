// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAIlIIl
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAIlllI
,
CAXI4DMAO0llI
,
CAXI4DMAI0llI
,
CAXI4DMAlOl1I
,
CAXI4DMAOIl1I
,
CAXI4DMAIIl1I
,
CAXI4DMAI1l1I
,
CAXI4DMAl1l1I
,
CAXI4DMAOO01I
,
CAXI4DMAlll1I
,
CAXI4DMAO0l1I
,
CAXI4DMAl100I
,
CAXI4DMAI0l1I
,
CAXI4DMAl0l1I
,
CAXI4DMAlIl1I
,
CAXI4DMAO1l1I
,
CAXI4DMAI1OOl
,
CAXI4DMAI1l1
,
CAXI4DMAlOlOl
,
CAXI4DMAIIllI
,
CAXI4DMAl1l1
,
CAXI4DMAOOOIl
,
strDscrptr
,
CAXI4DMAllllI
,
CAXI4DMAI1IlI
,
CAXI4DMAIIIIl
,
CAXI4DMAOIOIl
,
CAXI4DMAlOOIl
,
CAXI4DMAlIlOl
,
CAXI4DMAOllOl
,
CAXI4DMAlIOIl
,
CAXI4DMAO0IIl
,
CAXI4DMAI0IIl
,
CAXI4DMAlI0OI
,
CAXI4DMAII0OI
,
CAXI4DMAOIOOI
,
CAXI4DMAl11Ol
,
CAXI4DMAOI0Ol
,
CAXI4DMAIlOIl
,
CAXI4DMAl01Ol
)
;
parameter
NUM_INT_BDS
=
0
;
parameter
CAXI4DMAOIO1
=
5
;
parameter
NUM_PRI_LVLS
=
1
;
parameter
CAXI4DMAl0OI
=
23
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAIlllI
;
input
CAXI4DMAO0llI
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0llI
;
input
[
31
:
0
]
CAXI4DMAlOl1I
;
input
CAXI4DMAOIl1I
;
input
CAXI4DMAIIl1I
;
input
[
31
:
0
]
CAXI4DMAI1l1I
;
input
[
1
:
0
]
CAXI4DMAl1l1I
;
input
[
2
:
0
]
CAXI4DMAOO01I
;
input
[
2
:
0
]
CAXI4DMAlll1I
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAO0l1I
;
input
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAl100I
;
input
CAXI4DMAI0l1I
;
input
CAXI4DMAl0l1I
;
input
CAXI4DMAlIl1I
;
input
[
31
:
0
]
CAXI4DMAO1l1I
;
input
[
1
:
0
]
CAXI4DMAI1OOl
;
input
CAXI4DMAI1l1
;
input
CAXI4DMAlOlOl
;
input
CAXI4DMAIIllI
;
input
CAXI4DMAl1l1
;
output
CAXI4DMAOOOIl
;
output
strDscrptr
;
output
CAXI4DMAI1IlI
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO0IIl
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0IIl
;
output
[
31
:
0
]
CAXI4DMAlI0OI
;
output
CAXI4DMAII0OI
;
output
[
1
:
0
]
CAXI4DMAIIIIl
;
output
[
2
:
0
]
CAXI4DMAOIOIl
;
output
[
2
:
0
]
CAXI4DMAlOOIl
;
output
[
31
:
0
]
CAXI4DMAlIlOl
;
output
[
31
:
0
]
CAXI4DMAOllOl
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAlIOIl
;
output
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAllllI
;
output
CAXI4DMAOIOOI
;
output
CAXI4DMAl11Ol
;
output
CAXI4DMAOI0Ol
;
output
[
31
:
0
]
CAXI4DMAIlOIl
;
output
CAXI4DMAl01Ol
;
reg
[
1
:
0
]
CAXI4DMAIO10l
;
reg
[
31
:
0
]
CAXI4DMAII11l
;
reg
CAXI4DMAlI11l
;
reg
CAXI4DMAOl11l
;
reg
[
31
:
0
]
CAXI4DMAIl11l
;
reg
[
1
:
0
]
CAXI4DMAll11l
;
reg
[
2
:
0
]
CAXI4DMAO011l
;
reg
[
2
:
0
]
CAXI4DMAI011l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl011l
;
reg
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAO111l
;
reg
CAXI4DMAI111l
;
reg
CAXI4DMAl111l
;
reg
CAXI4DMAOOOO0
;
reg
[
31
:
0
]
CAXI4DMAIOOO0
;
reg
[
31
:
0
]
CAXI4DMAlOOO0
;
reg
CAXI4DMAOIOO0
;
reg
CAXI4DMAIIOO0
;
reg
[
31
:
0
]
CAXI4DMAlIOO0
;
reg
[
1
:
0
]
CAXI4DMAOlOO0
;
reg
[
2
:
0
]
CAXI4DMAIlOO0
;
reg
[
2
:
0
]
CAXI4DMAllOO0
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAO0OO0
;
reg
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAI0OO0
;
reg
CAXI4DMAl0OO0
;
reg
CAXI4DMAO1OO0
;
reg
CAXI4DMAI1OO0
;
reg
[
31
:
0
]
CAXI4DMAl1OO0
;
reg
[
1
:
0
]
CAXI4DMAO01Il
;
reg
CAXI4DMAl0O1l
;
reg
CAXI4DMAOOIO0
;
reg
CAXI4DMAIOIO0
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO10l
<=
2
'b
0
;
end
else
begin
case
(
{
CAXI4DMAIlllI
,
CAXI4DMAI1OOl
[
1
]
,
CAXI4DMAI1OOl
[
0
]
}
)
3
'b
000
,
3
'b
101
,
3
'b
110
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
;
end
3
'b
001
,
3
'b
010
,
3
'b
111
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
-
1
'b
1
;
end
3
'b
011
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
-
2
'b
10
;
end
3
'b
100
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
+
1
'b
1
;
end
endcase
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO01Il
[
1
:
0
]
<=
2
'b
0
;
end
else
begin
if
(
(
CAXI4DMAlOlOl
&
CAXI4DMAIIllI
)
||
(
CAXI4DMAO0llI
)
)
begin
CAXI4DMAO01Il
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
end
else
if
(
|
CAXI4DMAI1OOl
==
1
'b
1
)
begin
CAXI4DMAO01Il
[
CAXI4DMAI1l1
]
<=
1
'b
0
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0O1l
<=
1
'b
0
;
end
else
if
(
CAXI4DMAIlllI
)
begin
CAXI4DMAl0O1l
<=
~
CAXI4DMAl0O1l
;
end
end
assign
CAXI4DMAOOOIl
=
(
CAXI4DMAIO10l
!=
2
'b
0
)
?
(
CAXI4DMAI1l1
==
1
'b
1
)
?
CAXI4DMAO01Il
[
1
]
:
CAXI4DMAO01Il
[
0
]
:
1
'b
0
;
assign
CAXI4DMAl01Ol
=
(
CAXI4DMAIO10l
<
2
'b
10
)
?
1
'b
1
:
1
'b
0
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOOIO0
<=
1
'b
0
;
CAXI4DMAO0IIl
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAII11l
<=
32
'b
0
;
CAXI4DMAlI11l
<=
1
'b
0
;
CAXI4DMAOl11l
<=
1
'b
0
;
CAXI4DMAIl11l
<=
32
'b
0
;
CAXI4DMAll11l
<=
2
'b
0
;
CAXI4DMAO011l
<=
3
'b
0
;
CAXI4DMAI011l
<=
3
'b
0
;
CAXI4DMAl011l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAO111l
<=
{
NUM_PRI_LVLS
{
1
'b
0
}
}
;
CAXI4DMAI111l
<=
1
'b
0
;
CAXI4DMAl111l
<=
1
'b
0
;
CAXI4DMAOOOO0
<=
1
'b
0
;
CAXI4DMAIOOO0
<=
32
'b
0
;
end
else
begin
if
(
CAXI4DMAIlllI
&
!
CAXI4DMAl0O1l
)
begin
CAXI4DMAOOIO0
<=
CAXI4DMAO0llI
;
CAXI4DMAO0IIl
<=
CAXI4DMAI0llI
;
CAXI4DMAII11l
<=
CAXI4DMAlOl1I
;
CAXI4DMAlI11l
<=
CAXI4DMAOIl1I
;
CAXI4DMAOl11l
<=
CAXI4DMAIIl1I
;
CAXI4DMAIl11l
<=
CAXI4DMAI1l1I
;
CAXI4DMAll11l
<=
CAXI4DMAl1l1I
;
CAXI4DMAO011l
<=
CAXI4DMAOO01I
;
CAXI4DMAI011l
<=
CAXI4DMAlll1I
;
CAXI4DMAl011l
<=
CAXI4DMAO0l1I
;
CAXI4DMAO111l
<=
CAXI4DMAl100I
;
CAXI4DMAI111l
<=
CAXI4DMAI0l1I
;
CAXI4DMAl111l
<=
CAXI4DMAl0l1I
;
CAXI4DMAOOOO0
<=
CAXI4DMAlIl1I
;
CAXI4DMAIOOO0
<=
CAXI4DMAO1l1I
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIOIO0
<=
1
'b
0
;
CAXI4DMAI0IIl
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAlOOO0
<=
32
'b
0
;
CAXI4DMAOIOO0
<=
1
'b
0
;
CAXI4DMAIIOO0
<=
1
'b
0
;
CAXI4DMAlIOO0
<=
32
'b
0
;
CAXI4DMAOlOO0
<=
2
'b
0
;
CAXI4DMAIlOO0
<=
3
'b
0
;
CAXI4DMAllOO0
<=
3
'b
0
;
CAXI4DMAO0OO0
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAI0OO0
<=
{
NUM_PRI_LVLS
{
1
'b
0
}
}
;
CAXI4DMAl0OO0
<=
1
'b
0
;
CAXI4DMAO1OO0
<=
1
'b
0
;
CAXI4DMAI1OO0
<=
1
'b
0
;
CAXI4DMAl1OO0
<=
32
'b
0
;
end
else
begin
if
(
CAXI4DMAIlllI
&
CAXI4DMAl0O1l
)
begin
CAXI4DMAIOIO0
<=
CAXI4DMAO0llI
;
CAXI4DMAI0IIl
<=
CAXI4DMAI0llI
;
CAXI4DMAlOOO0
<=
CAXI4DMAlOl1I
;
CAXI4DMAOIOO0
<=
CAXI4DMAOIl1I
;
CAXI4DMAIIOO0
<=
CAXI4DMAIIl1I
;
CAXI4DMAlIOO0
<=
CAXI4DMAI1l1I
;
CAXI4DMAOlOO0
<=
CAXI4DMAl1l1I
;
CAXI4DMAIlOO0
<=
CAXI4DMAOO01I
;
CAXI4DMAllOO0
<=
CAXI4DMAlll1I
;
CAXI4DMAO0OO0
<=
CAXI4DMAO0l1I
;
CAXI4DMAI0OO0
<=
CAXI4DMAl100I
;
CAXI4DMAl0OO0
<=
CAXI4DMAI0l1I
;
CAXI4DMAO1OO0
<=
CAXI4DMAl0l1I
;
CAXI4DMAI1OO0
<=
CAXI4DMAlIl1I
;
CAXI4DMAl1OO0
<=
CAXI4DMAO1l1I
;
end
end
end
assign
strDscrptr
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAIOIO0
:
CAXI4DMAOOIO0
;
assign
CAXI4DMAIIIIl
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAOlOO0
:
CAXI4DMAll11l
;
assign
CAXI4DMAlI0OI
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAlOOO0
:
CAXI4DMAII11l
;
assign
CAXI4DMAII0OI
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAOIOO0
:
CAXI4DMAlI11l
;
assign
CAXI4DMAI1IlI
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAIIOO0
:
CAXI4DMAOl11l
;
assign
CAXI4DMAOIOIl
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAIlOO0
:
CAXI4DMAO011l
;
assign
CAXI4DMAlOOIl
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAllOO0
:
CAXI4DMAI011l
;
assign
CAXI4DMAlIlOl
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAlIOO0
:
CAXI4DMAIl11l
;
assign
CAXI4DMAlIOIl
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAO0OO0
:
CAXI4DMAl011l
;
assign
CAXI4DMAllllI
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAI0OO0
:
CAXI4DMAO111l
;
assign
CAXI4DMAOIOOI
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAl0OO0
:
CAXI4DMAI111l
;
assign
CAXI4DMAl11Ol
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAO1OO0
:
CAXI4DMAl111l
;
assign
CAXI4DMAOI0Ol
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAI1OO0
:
CAXI4DMAOOOO0
;
assign
CAXI4DMAIlOIl
=
(
CAXI4DMAI1l1
)
?
CAXI4DMAl1OO0
:
CAXI4DMAIOOO0
;
assign
CAXI4DMAOllOl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAlIOO0
:
CAXI4DMAIl11l
;
endmodule
