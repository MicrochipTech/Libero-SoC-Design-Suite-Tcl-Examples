// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAOOO1I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAO0I0I
,
CAXI4DMAlOO1I
,
CAXI4DMAl0I0I
,
CAXI4DMAO1I0I
,
CAXI4DMAI1I0I
,
CAXI4DMAOIO1I
,
CAXI4DMAIIO1I
,
CAXI4DMAl0IOI
,
CAXI4DMAl1I0I
,
CAXI4DMAOOl0I
,
CAXI4DMAIOl0I
,
CAXI4DMAlOl0I
,
CAXI4DMAOIl0I
,
CAXI4DMAIIl0I
,
CAXI4DMAlIl0I
,
CAXI4DMAllI0I
,
CAXI4DMAOll0I
,
CAXI4DMAIll0I
,
CAXI4DMAI1l0I
,
CAXI4DMAO010I
,
CAXI4DMAI010I
,
CAXI4DMAl1l0I
,
CAXI4DMAl0IlI
,
CAXI4DMAI1IlI
,
strDscrptr
,
CAXI4DMAlIO1I
,
intDscrptrNum
,
CAXI4DMAlI0OI
,
CAXI4DMAO1IOI
,
CAXI4DMAOlO1I
,
CAXI4DMAI0IOI
,
CAXI4DMAIlO1I
)
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl1OI
=
133
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAO0I0I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlOO1I
;
input
CAXI4DMAl0I0I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO1I0I
;
input
CAXI4DMAI1I0I
;
input
CAXI4DMAOIO1I
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAIIO1I
;
input
CAXI4DMAl0IOI
;
input
CAXI4DMAl1I0I
;
input
CAXI4DMAOOl0I
;
input
CAXI4DMAIOl0I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlOl0I
;
input
[
31
:
0
]
CAXI4DMAOIl0I
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAIIl0I
;
input
CAXI4DMAlIl0I
;
output
reg
CAXI4DMAllI0I
;
output
reg
CAXI4DMAOll0I
;
output
reg
CAXI4DMAIll0I
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI1l0I
;
output
reg
CAXI4DMAO010I
;
output
reg
CAXI4DMAI010I
;
output
reg
[
31
:
0
]
CAXI4DMAl1l0I
;
output
reg
CAXI4DMAl0IlI
;
output
reg
CAXI4DMAI1IlI
;
output
reg
strDscrptr
;
output
reg
CAXI4DMAlIO1I
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
intDscrptrNum
;
output
reg
[
31
:
0
]
CAXI4DMAlI0OI
;
output
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
output
reg
CAXI4DMAOlO1I
;
output
reg
CAXI4DMAI0IOI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIlO1I
;
localparam
[
1
:
0
]
CAXI4DMAI1lIl
=
2
'b
00
;
localparam
[
1
:
0
]
CAXI4DMAl1lIl
=
2
'b
01
;
localparam
[
1
:
0
]
CAXI4DMAOO0Il
=
2
'b
10
;
localparam
[
4
:
0
]
CAXI4DMAO1OII
=
5
'b
00001
;
localparam
[
4
:
0
]
CAXI4DMAIO0Il
=
5
'b
00010
;
localparam
[
4
:
0
]
CAXI4DMAlO0Il
=
5
'b
00100
;
localparam
[
4
:
0
]
CAXI4DMAOI0Il
=
5
'b
01000
;
localparam
[
4
:
0
]
CAXI4DMAII0Il
=
5
'b
10000
;
wire
[
2
:
0
]
CAXI4DMAlI0Il
;
wire
[
2
:
0
]
CAXI4DMAIlO0I
;
reg
CAXI4DMAlI11I
;
wire
[
1
:
0
]
CAXI4DMAOl0Il
;
reg
CAXI4DMAIl0Il
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAll0Il
;
reg
CAXI4DMAO00Il
;
reg
CAXI4DMAI00Il
;
reg
[
31
:
0
]
CAXI4DMAl00Il
;
reg
CAXI4DMAO10Il
;
reg
[
4
:
0
]
CAXI4DMAl10OI
;
reg
[
4
:
0
]
CAXI4DMAOO1OI
;
CAXI4DMAOI11I
#
(
.CAXI4DMAIl1lI
(
3
)
)
CAXI4DMAI10Il
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
CAXI4DMAlI0Il
)
,
.CAXI4DMAlI11I
(
CAXI4DMAlI11I
)
,
.CAXI4DMAOl11I
(
)
,
.CAXI4DMAIlO0I
(
CAXI4DMAIlO0I
)
)
;
assign
CAXI4DMAlI0Il
=
{
CAXI4DMAl1I0I
,
CAXI4DMAl0I0I
,
CAXI4DMAO0I0I
}
;
assign
CAXI4DMAOl0Il
=
(
CAXI4DMAIlO0I
==
3
'b
010
)
?
CAXI4DMAl1lIl
:
(
CAXI4DMAIlO0I
==
3
'b
100
)
?
CAXI4DMAOO0Il
:
CAXI4DMAI1lIl
;
assign
CAXI4DMAIlO1I
=
(
CAXI4DMAOl0Il
[
0
]
)
?
CAXI4DMAO1I0I
:
CAXI4DMAlOO1I
;
always
@
(
*
)
begin
case
(
CAXI4DMAOl0Il
)
CAXI4DMAI1lIl
:
begin
CAXI4DMAO10Il
<=
CAXI4DMAOIO1I
;
CAXI4DMAI1IlI
<=
1
'b
0
;
strDscrptr
<=
1
'b
0
;
CAXI4DMAlIO1I
<=
1
'b
0
;
intDscrptrNum
<=
CAXI4DMAIlO1I
;
CAXI4DMAlI0OI
<=
32
'b
0
;
CAXI4DMAO1IOI
<=
CAXI4DMAIIO1I
;
end
CAXI4DMAl1lIl
:
begin
CAXI4DMAO10Il
<=
CAXI4DMAOIO1I
;
CAXI4DMAI1IlI
<=
1
'b
0
;
strDscrptr
<=
1
'b
0
;
CAXI4DMAlIO1I
<=
1
'b
0
;
intDscrptrNum
<=
CAXI4DMAIlO1I
;
CAXI4DMAlI0OI
<=
32
'b
0
;
CAXI4DMAO1IOI
<=
CAXI4DMAIIO1I
;
end
CAXI4DMAOO0Il
:
begin
CAXI4DMAO10Il
<=
CAXI4DMAlIl0I
;
CAXI4DMAI1IlI
<=
CAXI4DMAOOl0I
;
strDscrptr
<=
CAXI4DMAIOl0I
;
CAXI4DMAlIO1I
<=
1
'b
1
;
intDscrptrNum
<=
CAXI4DMAlOl0I
;
CAXI4DMAlI0OI
<=
CAXI4DMAOIl0I
;
CAXI4DMAO1IOI
<=
CAXI4DMAIIl0I
;
end
default
:
begin
CAXI4DMAO10Il
<=
1
'b
0
;
CAXI4DMAI1IlI
<=
1
'b
0
;
strDscrptr
<=
1
'b
0
;
CAXI4DMAlIO1I
<=
1
'b
0
;
intDscrptrNum
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAlI0OI
<=
32
'b
0
;
CAXI4DMAO1IOI
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAI0IOI
<=
1
'b
0
;
CAXI4DMAllI0I
<=
1
'b
0
;
CAXI4DMAOll0I
<=
1
'b
0
;
CAXI4DMAOlO1I
<=
1
'b
0
;
CAXI4DMAl0IlI
<=
1
'b
0
;
CAXI4DMAlI11I
<=
1
'b
0
;
CAXI4DMAIl0Il
<=
1
'b
0
;
CAXI4DMAll0Il
<=
CAXI4DMAI1l0I
;
CAXI4DMAO00Il
<=
CAXI4DMAO010I
;
CAXI4DMAI00Il
<=
CAXI4DMAI010I
;
CAXI4DMAl00Il
<=
CAXI4DMAl1l0I
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
|
CAXI4DMAIlO0I
[
2
:
0
]
)
begin
if
(
|
CAXI4DMAIlO0I
[
1
:
0
]
)
begin
CAXI4DMAI0IOI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO0Il
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOI0Il
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAIO0Il
:
begin
if
(
CAXI4DMAl0IOI
)
begin
if
(
CAXI4DMAO10Il
)
begin
CAXI4DMAl0IlI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAII0Il
;
end
else
begin
CAXI4DMAIl0Il
<=
1
'b
1
;
CAXI4DMAll0Il
<=
intDscrptrNum
;
CAXI4DMAO00Il
<=
1
'b
0
;
CAXI4DMAI00Il
<=
1
'b
0
;
CAXI4DMAl00Il
<=
32
'b
0
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO0Il
;
end
if
(
CAXI4DMAIlO0I
[
0
]
)
begin
CAXI4DMAllI0I
<=
1
'b
1
;
end
else
if
(
CAXI4DMAIlO0I
[
1
]
)
begin
CAXI4DMAOll0I
<=
1
'b
1
;
end
end
else
begin
CAXI4DMAI0IOI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO0Il
;
end
end
CAXI4DMAOI0Il
:
begin
CAXI4DMAOlO1I
<=
1
'b
1
;
if
(
CAXI4DMAO10Il
)
begin
CAXI4DMAl0IlI
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAII0Il
;
end
else
begin
CAXI4DMAIl0Il
<=
1
'b
1
;
CAXI4DMAll0Il
<=
intDscrptrNum
;
CAXI4DMAO00Il
<=
CAXI4DMAlIO1I
;
CAXI4DMAI00Il
<=
strDscrptr
;
CAXI4DMAl00Il
<=
CAXI4DMAlI0OI
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO0Il
;
end
end
CAXI4DMAlO0Il
:
begin
if
(
CAXI4DMAI1I0I
)
begin
CAXI4DMAlI11I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAIl0Il
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO0Il
;
end
end
CAXI4DMAII0Il
:
begin
CAXI4DMAlI11I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIll0I
<=
1
'b
0
;
end
else
begin
CAXI4DMAIll0I
<=
CAXI4DMAIl0Il
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1l0I
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAI1l0I
<=
CAXI4DMAll0Il
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl1l0I
<=
32
'b
0
;
end
else
begin
CAXI4DMAl1l0I
<=
CAXI4DMAl00Il
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO010I
<=
1
'b
0
;
end
else
begin
CAXI4DMAO010I
<=
CAXI4DMAO00Il
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI010I
<=
1
'b
0
;
end
else
begin
CAXI4DMAI010I
<=
CAXI4DMAI00Il
;
end
end
endmodule
