// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAIOIIl
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAIlllI
,
CAXI4DMAOll0I
,
CAXI4DMAOl0
,
CAXI4DMAlI1Ol
,
CAXI4DMAl00Ol
,
CAXI4DMAlOlOl
,
CAXI4DMAOIlOl
,
CAXI4DMAOIIIl
,
CAXI4DMAl01Ol
,
CAXI4DMAIIIIl
,
CAXI4DMAlIIIl
,
CAXI4DMAIOOOl
,
CAXI4DMAOlOIl
,
CAXI4DMAOIOOI
,
CAXI4DMAl11Ol
,
CAXI4DMAII0OI
,
CAXI4DMAIOOIl
,
CAXI4DMAOOlOl
,
CAXI4DMAIOlOl
,
CAXI4DMAOIOOl
,
CAXI4DMAIIOOl
,
CAXI4DMAOlIIl
,
CAXI4DMAl1l1
,
CAXI4DMAlOllI
,
strDscrptr
,
CAXI4DMAIIllI
,
CAXI4DMAl1IlI
,
CAXI4DMAOOllI
,
CAXI4DMAIOllI
,
CAXI4DMAl0I0I
,
intDscrptrNum
)
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl0OI
=
4
;
parameter
CAXI4DMAO1OI
=
13
;
parameter
AXI4_STREAM_IF
=
0
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAIlllI
;
input
CAXI4DMAOll0I
;
input
CAXI4DMAOl0
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI1Ol
;
input
CAXI4DMAl00Ol
;
input
CAXI4DMAlOlOl
;
input
CAXI4DMAOIlOl
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAOIIIl
;
input
CAXI4DMAl01Ol
;
input
[
1
:
0
]
CAXI4DMAIIIIl
;
input
[
31
:
0
]
CAXI4DMAlIIIl
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIOOOl
;
input
CAXI4DMAOlOIl
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOIOOl
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIIOOl
;
input
CAXI4DMAOIOOI
;
input
CAXI4DMAl11Ol
;
input
CAXI4DMAII0OI
;
input
[
1
:
0
]
CAXI4DMAIOOIl
;
input
[
31
:
0
]
CAXI4DMAOOlOl
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIOlOl
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOlIIl
;
input
CAXI4DMAl1l1
;
output
CAXI4DMAlOllI
;
output
strDscrptr
;
output
CAXI4DMAIIllI
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl1IlI
;
output
[
31
:
0
]
CAXI4DMAOOllI
;
output
[
31
:
0
]
CAXI4DMAIOllI
;
output
CAXI4DMAl0I0I
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
intDscrptrNum
;
reg
[
2
:
0
]
CAXI4DMAl10OI
;
reg
[
2
:
0
]
CAXI4DMAOO1OI
;
reg
CAXI4DMAIlI1l
;
reg
CAXI4DMAllI1l
;
reg
CAXI4DMAIO00l
;
reg
CAXI4DMAlO00l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAO0I1l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAI0I1l
;
reg
[
31
:
0
]
CAXI4DMAl0I1l
;
reg
[
31
:
0
]
CAXI4DMAO1I1l
;
reg
[
31
:
0
]
CAXI4DMAI1I1l
;
reg
[
31
:
0
]
CAXI4DMAl1I1l
;
reg
CAXI4DMAOOl1l
;
reg
CAXI4DMAIOl1l
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl01Il
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO11Il
;
reg
CAXI4DMAlOl1l
;
reg
CAXI4DMAOIl1l
;
localparam
[
2
:
0
]
CAXI4DMAO1OII
=
3
'b
001
;
localparam
[
2
:
0
]
CAXI4DMAIIl1l
=
3
'b
010
;
localparam
[
2
:
0
]
CAXI4DMAlIl1l
=
3
'b
100
;
localparam
[
1
:
0
]
CAXI4DMAOll1l
=
2
'b
01
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAIOl1l
<=
1
'b
0
;
CAXI4DMAO11Il
<=
CAXI4DMAl01Il
;
CAXI4DMAlO00l
<=
CAXI4DMAIO00l
;
CAXI4DMAllI1l
<=
1
'b
0
;
CAXI4DMAI0I1l
<=
CAXI4DMAO0I1l
;
CAXI4DMAO1I1l
<=
CAXI4DMAl0I1l
;
CAXI4DMAl1I1l
<=
CAXI4DMAI1I1l
;
CAXI4DMAOIl1l
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAIlllI
)
begin
if
(
CAXI4DMAl01Ol
&
CAXI4DMAOlOIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIIl1l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAIIl1l
:
begin
if
(
CAXI4DMAlOlOl
)
begin
CAXI4DMAllI1l
<=
1
'b
1
;
CAXI4DMAOIl1l
<=
1
'b
0
;
CAXI4DMAlO00l
<=
CAXI4DMAOIlOl
;
if
(
CAXI4DMAIOOIl
==
2
'b
00
)
begin
CAXI4DMAI0I1l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAO1I1l
<=
CAXI4DMAOOlOl
;
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
if
(
CAXI4DMAOIOOI
)
begin
if
(
!
CAXI4DMAl11Ol
)
begin
CAXI4DMAIOl1l
<=
1
'b
1
;
CAXI4DMAO11Il
<=
CAXI4DMAOlIIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAlIl1l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
if
(
CAXI4DMAII0OI
)
begin
if
(
CAXI4DMAOIlOl
)
begin
CAXI4DMAI0I1l
<=
CAXI4DMAIOlOl
-
CAXI4DMAOIIIl
;
if
(
CAXI4DMAIOOIl
==
CAXI4DMAOll1l
)
begin
CAXI4DMAO1I1l
<=
CAXI4DMAOOlOl
+
CAXI4DMAOIIIl
;
end
else
begin
CAXI4DMAO1I1l
<=
CAXI4DMAOOlOl
;
end
if
(
CAXI4DMAIIIIl
==
CAXI4DMAOll1l
)
begin
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
+
CAXI4DMAOIIIl
;
end
else
begin
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
end
if
(
CAXI4DMAIOlOl
==
{
{
(
CAXI4DMAl0OI
-
CAXI4DMAO1OI
)
{
1
'b
0
}
}
,
CAXI4DMAOIIIl
}
)
begin
if
(
CAXI4DMAOIOOI
)
begin
if
(
!
CAXI4DMAl11Ol
)
begin
CAXI4DMAIOl1l
<=
1
'b
1
;
CAXI4DMAO11Il
<=
CAXI4DMAOlIIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAlIl1l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAI0I1l
<=
CAXI4DMAIOlOl
;
CAXI4DMAO1I1l
<=
CAXI4DMAOOlOl
;
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAI0I1l
<=
CAXI4DMAIOlOl
-
CAXI4DMAOIIIl
;
if
(
CAXI4DMAIOOIl
==
CAXI4DMAOll1l
)
begin
CAXI4DMAO1I1l
<=
CAXI4DMAOOlOl
+
CAXI4DMAOIIIl
;
end
else
begin
CAXI4DMAO1I1l
<=
CAXI4DMAOOlOl
;
end
if
(
CAXI4DMAIIIIl
==
CAXI4DMAOll1l
)
begin
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
+
CAXI4DMAOIIIl
;
end
else
begin
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
end
if
(
CAXI4DMAIOlOl
==
{
{
(
CAXI4DMAl0OI
-
CAXI4DMAO1OI
)
{
1
'b
0
}
}
,
CAXI4DMAOIIIl
}
)
begin
if
(
CAXI4DMAOIOOI
)
begin
if
(
!
CAXI4DMAl11Ol
)
begin
CAXI4DMAIOl1l
<=
1
'b
1
;
CAXI4DMAO11Il
<=
CAXI4DMAOlIIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAlIl1l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
end
else
if
(
(
CAXI4DMAOl0
==
1
'b
1
)
&&
(
AXI4_STREAM_IF
==
1
)
)
begin
CAXI4DMAllI1l
<=
1
'b
1
;
CAXI4DMAOIl1l
<=
1
'b
1
;
CAXI4DMAlO00l
<=
1
'b
1
;
CAXI4DMAI0I1l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
if
(
CAXI4DMAIIIIl
==
CAXI4DMAOll1l
)
begin
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
+
CAXI4DMAlI1Ol
;
end
else
begin
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
end
end
else
if
(
(
CAXI4DMAl00Ol
==
1
'b
1
)
&&
(
AXI4_STREAM_IF
==
1
)
)
begin
CAXI4DMAllI1l
<=
1
'b
1
;
CAXI4DMAOIl1l
<=
1
'b
1
;
CAXI4DMAlO00l
<=
1
'b
0
;
CAXI4DMAI0I1l
<=
CAXI4DMAIOOOl
;
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
CAXI4DMAl1I1l
<=
CAXI4DMAlIIIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIIl1l
;
end
end
CAXI4DMAlIl1l
:
begin
if
(
CAXI4DMAOll0I
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAIOl1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlIl1l
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIlI1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAIlI1l
<=
CAXI4DMAllI1l
;
end
end
assign
CAXI4DMAlOllI
=
CAXI4DMAIlI1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO00l
<=
1
'b
0
;
end
else
begin
CAXI4DMAIO00l
<=
CAXI4DMAlO00l
;
end
end
assign
CAXI4DMAIIllI
=
CAXI4DMAIO00l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO0I1l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAO0I1l
<=
CAXI4DMAI0I1l
;
end
end
assign
CAXI4DMAl1IlI
=
CAXI4DMAO0I1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0I1l
<=
32
'b
0
;
end
else
begin
CAXI4DMAl0I1l
<=
CAXI4DMAO1I1l
;
end
end
assign
CAXI4DMAOOllI
=
CAXI4DMAl0I1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1I1l
<=
32
'b
0
;
end
else
begin
CAXI4DMAI1I1l
<=
CAXI4DMAl1I1l
;
end
end
assign
CAXI4DMAIOllI
=
CAXI4DMAI1I1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOOl1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAOOl1l
<=
CAXI4DMAIOl1l
;
end
end
assign
CAXI4DMAl0I0I
=
CAXI4DMAOOl1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl01Il
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAl01Il
<=
CAXI4DMAO11Il
;
end
end
assign
intDscrptrNum
=
CAXI4DMAl01Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlOl1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAlOl1l
<=
CAXI4DMAOIl1l
;
end
end
assign
strDscrptr
=
CAXI4DMAlOl1l
;
endmodule
