// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAl1I1I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAIOl1I
,
CAXI4DMAO0llI
,
CAXI4DMAI0llI
,
CAXI4DMAlOl1I
,
CAXI4DMAOIl1I
,
CAXI4DMAl100I
,
CAXI4DMAIIl1I
,
CAXI4DMAlIl1I
,
CAXI4DMAOll1I
,
CAXI4DMAIll1I
,
CAXI4DMAlll1I
,
CAXI4DMAO0l1I
,
CAXI4DMAI0l1I
,
CAXI4DMAl0l1I
,
CAXI4DMAO1l1I
,
CAXI4DMAI1l1I
,
CAXI4DMAl1l1I
,
CAXI4DMAOO01I
,
CAXI4DMAII10I
,
CAXI4DMAIO01I
,
CAXI4DMAlO01I
,
CAXI4DMAOI01I
,
CAXI4DMAII01I
,
CAXI4DMAlO0
,
CAXI4DMAOI0
,
CAXI4DMAl011
,
CAXI4DMAO111
,
CAXI4DMAOl0
,
CAXI4DMAIl0
,
CAXI4DMAll0
,
CAXI4DMAO00
,
CAXI4DMAI00
,
CAXI4DMAlI01I
,
CAXI4DMAOl01I
,
CAXI4DMAlI10I
,
CAXI4DMAll00I
,
CAXI4DMAO000I
,
CAXI4DMAIl01I
,
CAXI4DMAlOllI
,
CAXI4DMAOIllI
,
CAXI4DMAIIllI
,
CAXI4DMAl1IlI
,
CAXI4DMAOOllI
,
CAXI4DMAIOllI
,
CAXI4DMAIO0lI
,
CAXI4DMAOlllI
,
CAXI4DMAOO10I
,
CAXI4DMAlIlOI
,
CAXI4DMAOllOI
,
CAXI4DMAIllOI
,
CAXI4DMAll01I
,
CAXI4DMAO001I
,
CAXI4DMAI001I
,
CAXI4DMAl001I
,
CAXI4DMAI1l1
,
CAXI4DMAl1l1
,
CAXI4DMAOI
,
CAXI4DMAII
,
CAXI4DMAlI
,
CAXI4DMAOl
,
CAXI4DMAll
,
CAXI4DMAO101I
,
CAXI4DMAO0
,
CAXI4DMAI0
,
CAXI4DMAl0
,
CAXI4DMAOIlOI
,
CAXI4DMAI1
,
CAXI4DMAI101I
,
CAXI4DMAOOI
,
CAXI4DMAIOI
,
CAXI4DMAlOI
,
CAXI4DMAOII
,
CAXI4DMAIII
,
CAXI4DMAlII
,
CAXI4DMAOlI
,
CAXI4DMAI0O1I
,
CAXI4DMAl0O1I
,
CAXI4DMAO1O1I
,
CAXI4DMAlOl0I
,
CAXI4DMAOIl0I
,
CAXI4DMAO1I
,
CAXI4DMAl0I0I
,
CAXI4DMAl0l0I
,
CAXI4DMAOl1l
,
CAXI4DMAIl1l
)
;
parameter
AXI4_STREAM_IF
=
0
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl0OI
=
23
;
parameter
CAXI4DMAO1OI
=
12
;
parameter
NUM_PRI_LVLS
=
1
;
parameter
CAXI4DMAI1OI
=
0
;
parameter
PRI_0_NUM_OF_BEATS
=
0
;
parameter
PRI_1_NUM_OF_BEATS
=
0
;
parameter
PRI_2_NUM_OF_BEATS
=
0
;
parameter
PRI_3_NUM_OF_BEATS
=
0
;
parameter
PRI_4_NUM_OF_BEATS
=
0
;
parameter
PRI_5_NUM_OF_BEATS
=
0
;
parameter
PRI_6_NUM_OF_BEATS
=
0
;
parameter
PRI_7_NUM_OF_BEATS
=
0
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAIOl1I
;
input
CAXI4DMAO0llI
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0llI
;
input
[
31
:
0
]
CAXI4DMAlOl1I
;
input
CAXI4DMAOIl1I
;
input
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAl100I
;
input
CAXI4DMAIIl1I
;
input
CAXI4DMAlIl1I
;
input
[
31
:
0
]
CAXI4DMAOll1I
;
input
[
1
:
0
]
CAXI4DMAIll1I
;
input
[
2
:
0
]
CAXI4DMAlll1I
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAO0l1I
;
input
CAXI4DMAI0l1I
;
input
CAXI4DMAl0l1I
;
input
[
31
:
0
]
CAXI4DMAO1l1I
;
input
[
31
:
0
]
CAXI4DMAI1l1I
;
input
[
1
:
0
]
CAXI4DMAl1l1I
;
input
[
2
:
0
]
CAXI4DMAOO01I
;
input
CAXI4DMAII10I
;
input
CAXI4DMAIO01I
;
input
CAXI4DMAlO01I
;
input
CAXI4DMAOI01I
;
input
CAXI4DMAII01I
;
input
CAXI4DMAlO0
;
input
CAXI4DMAOI0
;
input
CAXI4DMAl011
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAO111
;
input
CAXI4DMAOl0
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIl0
;
input
CAXI4DMAll0
;
input
CAXI4DMAO00
;
input
CAXI4DMAI00
;
input
CAXI4DMAlI01I
;
input
CAXI4DMAOl01I
;
input
CAXI4DMAlI10I
;
input
CAXI4DMAll00I
;
input
CAXI4DMAO000I
;
input
CAXI4DMAIl01I
;
output
CAXI4DMAlOllI
;
output
CAXI4DMAOIllI
;
output
CAXI4DMAIIllI
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl1IlI
;
output
[
31
:
0
]
CAXI4DMAOOllI
;
output
[
31
:
0
]
CAXI4DMAIOllI
;
output
CAXI4DMAIO0lI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOlllI
;
output
CAXI4DMAOO10I
;
output
CAXI4DMAlIlOI
;
output
CAXI4DMAOllOI
;
output
CAXI4DMAIllOI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAll01I
;
output
CAXI4DMAO001I
;
output
[
31
:
0
]
CAXI4DMAI001I
;
output
CAXI4DMAl001I
;
output
CAXI4DMAI1l1
;
output
CAXI4DMAl1l1
;
output
CAXI4DMAOI
;
output
CAXI4DMAII
;
output
[
1
:
0
]
CAXI4DMAlI
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOl
;
output
[
2
:
0
]
CAXI4DMAll
;
output
[
31
:
0
]
CAXI4DMAO101I
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAO0
;
output
CAXI4DMAI0
;
output
[
1
:
0
]
CAXI4DMAl0
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOIlOI
;
output
[
2
:
0
]
CAXI4DMAI1
;
output
[
31
:
0
]
CAXI4DMAI101I
;
output
[
2
:
0
]
CAXI4DMAOOI
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAIOI
;
output
CAXI4DMAlOI
;
output
[
31
:
0
]
CAXI4DMAOII
;
output
CAXI4DMAIII
;
output
[
31
:
0
]
CAXI4DMAlII
;
output
[
1
:
0
]
CAXI4DMAOlI
;
output
CAXI4DMAI0O1I
;
output
CAXI4DMAl0O1I
;
output
CAXI4DMAO1O1I
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlOl0I
;
output
[
31
:
0
]
CAXI4DMAOIl0I
;
output
[
7
:
0
]
CAXI4DMAO1I
;
output
CAXI4DMAl0I0I
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl0l0I
;
output
CAXI4DMAOl1l
;
output
CAXI4DMAIl1l
;
wire
[
31
:
0
]
CAXI4DMAIl11I
;
wire
[
31
:
0
]
CAXI4DMAll11I
;
wire
CAXI4DMAO011I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI011I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl011I
;
wire
[
31
:
0
]
CAXI4DMAO111I
;
wire
CAXI4DMAI111I
;
wire
CAXI4DMAl111I
;
wire
CAXI4DMAOOOOl
;
wire
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIOOOl
;
wire
CAXI4DMAlOOOl
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOIOOl
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIIOOl
;
wire
[
31
:
0
]
CAXI4DMAlIOOl
;
wire
CAXI4DMAOlOOl
;
wire
CAXI4DMAIlOOl
;
wire
CAXI4DMAllOOl
;
wire
CAXI4DMAO0OOl
;
wire
CAXI4DMAI0OOl
;
wire
CAXI4DMAl0OOl
;
wire
CAXI4DMAO1OOl
;
wire
[
1
:
0
]
CAXI4DMAI1OOl
;
wire
[
1
:
0
]
CAXI4DMAl1OOl
;
wire
CAXI4DMAOOIOl
;
wire
CAXI4DMAIOIOl
;
wire
CAXI4DMAlOIOl
;
wire
CAXI4DMAOIIOl
;
wire
CAXI4DMAIIIOl
;
wire
CAXI4DMAlIIOl
;
wire
CAXI4DMAOlIOl
;
wire
[
31
:
0
]
CAXI4DMAIlIOl
;
wire
CAXI4DMAllIOl
;
wire
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAO0IOl
;
wire
CAXI4DMAI0IOl
;
wire
CAXI4DMAl0IOl
;
wire
[
1
:
0
]
CAXI4DMAO1IOl
;
wire
[
2
:
0
]
CAXI4DMAI1IOl
;
wire
[
2
:
0
]
CAXI4DMAl1IOl
;
wire
[
31
:
0
]
CAXI4DMAOOlOl
;
wire
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIOlOl
;
wire
CAXI4DMAlOlOl
;
wire
CAXI4DMAOIlOl
;
wire
[
1
:
0
]
CAXI4DMAIIlOl
;
wire
[
31
:
0
]
CAXI4DMAlIlOl
;
wire
[
31
:
0
]
CAXI4DMAOllOl
;
wire
CAXI4DMAIllOl
;
wire
[
2
:
0
]
CAXI4DMAlllOl
;
wire
[
2
:
0
]
CAXI4DMAO0lOl
;
wire
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAI0lOl
;
wire
CAXI4DMAl0lOl
;
wire
CAXI4DMAO1lOl
;
wire
[
7
:
0
]
CAXI4DMAI1lOl
;
wire
CAXI4DMAl1lOl
;
wire
CAXI4DMAOO0Ol
;
wire
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIO0Ol
;
wire
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlO0Ol
;
wire
CAXI4DMAOI0Ol
;
reg
[
1
:
0
]
CAXI4DMAII0Ol
;
reg
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI0Ol
[
0
:
1
]
;
reg
CAXI4DMAl10OI
;
reg
CAXI4DMAOO1OI
;
reg
CAXI4DMAOl0Ol
;
wire
[
31
:
0
]
CAXI4DMAIl0Ol
;
wire
CAXI4DMAll0Ol
;
wire
CAXI4DMAO00Ol
;
wire
CAXI4DMAI00Ol
;
wire
CAXI4DMAl00Ol
;
wire
CAXI4DMAO10Ol
;
wire
CAXI4DMAI10Ol
;
wire
CAXI4DMAl10Ol
;
wire
CAXI4DMAOO1Ol
;
localparam
CAXI4DMAO1OII
=
1
'b
0
;
localparam
CAXI4DMAIO1Ol
=
1
'b
1
;
assign
CAXI4DMAOIl0I
=
(
CAXI4DMAO1O1I
)
?
CAXI4DMAIl11I
:
CAXI4DMAll11I
;
assign
CAXI4DMAI1lOl
=
{
1
'b
1
,
1
'b
0
,
1
'b
0
,
CAXI4DMAOI0Ol
,
CAXI4DMAO1lOl
,
CAXI4DMAl0lOl
,
CAXI4DMAlllOl
[
2
:
1
]
}
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAIOl1I
&
CAXI4DMAlOOOl
&
CAXI4DMAO011I
)
begin
CAXI4DMAOl0Ol
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO1Ol
;
end
else
begin
CAXI4DMAOl0Ol
<=
1
'b
0
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAIO1Ol
:
begin
CAXI4DMAOl0Ol
<=
1
'b
0
;
if
(
CAXI4DMAlOllI
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIO1Ol
;
end
end
endcase
end
CAXI4DMAlO1Ol
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAO1OI
(
CAXI4DMAO1OI
)
)
CAXI4DMAOI1Ol
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO011I
(
CAXI4DMAO011I
)
,
.CAXI4DMAI011I
(
CAXI4DMAI011I
)
,
.CAXI4DMAl011I
(
CAXI4DMAl011I
)
,
.CAXI4DMAO111I
(
CAXI4DMAO111I
)
,
.CAXI4DMAI111I
(
CAXI4DMAI111I
)
,
.CAXI4DMAII1Ol
(
CAXI4DMAIl0Ol
)
,
.CAXI4DMAIOOOl
(
CAXI4DMAIOOOl
)
,
.CAXI4DMAI1lOl
(
CAXI4DMAI1lOl
)
,
.CAXI4DMAOI0Ol
(
CAXI4DMAOI0Ol
)
,
.CAXI4DMAl0lOl
(
CAXI4DMAl0lOl
)
,
.CAXI4DMAO1lOl
(
CAXI4DMAO1lOl
)
,
.CAXI4DMAIIlOl
(
CAXI4DMAIIlOl
)
,
.CAXI4DMAlOOOl
(
CAXI4DMAlOOOl
)
,
.CAXI4DMAI0IOl
(
CAXI4DMAI0IOl
)
,
.CAXI4DMAl111I
(
CAXI4DMAl111I
)
,
.CAXI4DMAOOOOl
(
CAXI4DMAOOOOl
)
,
.CAXI4DMAOIOOl
(
CAXI4DMAOIOOl
)
,
.CAXI4DMAIIOOl
(
CAXI4DMAIIOOl
)
,
.CAXI4DMAlIOOl
(
CAXI4DMAlIOOl
)
,
.CAXI4DMAIOlOl
(
CAXI4DMAIOlOl
)
,
.CAXI4DMAlI0
(
CAXI4DMAIO0Ol
)
,
.CAXI4DMAOlOOl
(
CAXI4DMAOlOOl
)
,
.CAXI4DMAIlOOl
(
CAXI4DMAIlOOl
)
,
.CAXI4DMAllOOl
(
CAXI4DMAllOOl
)
,
.CAXI4DMAO0OOl
(
CAXI4DMAO0OOl
)
,
.CAXI4DMAlI1Ol
(
CAXI4DMAlO0Ol
)
,
.CAXI4DMAI00
(
CAXI4DMAI00
)
,
.CAXI4DMAI10Ol
(
CAXI4DMAI10Ol
)
,
.CAXI4DMAl00Ol
(
CAXI4DMAl00Ol
)
,
.CAXI4DMAI0OOl
(
CAXI4DMAI0OOl
)
,
.CAXI4DMAl0OOl
(
CAXI4DMAl0OOl
)
,
.CAXI4DMAO1OOl
(
CAXI4DMAO1OOl
)
,
.CAXI4DMAO10Ol
(
CAXI4DMAO10Ol
)
,
.CAXI4DMAI1I1I
(
CAXI4DMAII10I
)
,
.CAXI4DMAOII1I
(
CAXI4DMAOl01I
)
,
.CAXI4DMAIII1I
(
CAXI4DMAlI10I
)
,
.CAXI4DMAIO0lI
(
CAXI4DMAIO0lI
)
,
.CAXI4DMAOlllI
(
CAXI4DMAOlllI
)
,
.CAXI4DMAI1OOl
(
CAXI4DMAI1OOl
)
,
.CAXI4DMAl1OOl
(
CAXI4DMAl1OOl
)
,
.CAXI4DMAOO10I
(
CAXI4DMAOO10I
)
,
.CAXI4DMAlIlOI
(
CAXI4DMAlIlOI
)
,
.CAXI4DMAOllOI
(
CAXI4DMAOllOI
)
,
.CAXI4DMAIllOI
(
CAXI4DMAIllOI
)
,
.CAXI4DMAI1l0I
(
CAXI4DMAll01I
)
,
.CAXI4DMAO010I
(
CAXI4DMAO001I
)
,
.CAXI4DMAl1l0I
(
CAXI4DMAI001I
)
,
.CAXI4DMAI010I
(
CAXI4DMAl001I
)
,
.CAXI4DMAOOIOl
(
CAXI4DMAOOIOl
)
,
.CAXI4DMAIOIOl
(
CAXI4DMAIOIOl
)
,
.CAXI4DMAlOIOl
(
CAXI4DMAlOIOl
)
,
.CAXI4DMAOIIOl
(
CAXI4DMAOIIOl
)
,
.CAXI4DMAIII
(
CAXI4DMAIII
)
,
.CAXI4DMAlII
(
CAXI4DMAlII
)
,
.CAXI4DMAOlI
(
CAXI4DMAOlI
)
,
.CAXI4DMAOO1Ol
(
CAXI4DMAOO1Ol
)
,
.CAXI4DMAIIIOl
(
CAXI4DMAIIIOl
)
,
.CAXI4DMAlIIOl
(
CAXI4DMAlIIOl
)
,
.CAXI4DMAOlIOl
(
CAXI4DMAOlIOl
)
,
.CAXI4DMAl10Ol
(
CAXI4DMAl10Ol
)
,
.CAXI4DMAI1l1
(
CAXI4DMAI1l1
)
,
.CAXI4DMAl1l1
(
CAXI4DMAl1l1
)
,
.CAXI4DMAOl1Ol
(
CAXI4DMAI0O1I
)
,
.CAXI4DMAl0I
(
CAXI4DMAl0O1I
)
,
.CAXI4DMAIl1Ol
(
CAXI4DMAlOl0I
)
,
.CAXI4DMAll1Ol
(
CAXI4DMAll11I
)
,
.CAXI4DMAO1I
(
CAXI4DMAO1I
)
,
.CAXI4DMAl1lOl
(
CAXI4DMAl1lOl
)
,
.CAXI4DMAOl1l
(
CAXI4DMAOl1l
)
,
.CAXI4DMAIl1l
(
CAXI4DMAIl1l
)
)
;
CAXI4DMAO01Ol
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.NUM_PRI_LVLS
(
NUM_PRI_LVLS
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
)
CAXI4DMAI01Ol
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAIlllI
(
CAXI4DMAOl0Ol
&
!
CAXI4DMAO0llI
)
,
.CAXI4DMAI0llI
(
CAXI4DMAI0llI
)
,
.CAXI4DMAlOl1I
(
CAXI4DMAlOl1I
)
,
.CAXI4DMAOIl1I
(
CAXI4DMAOIl1I
)
,
.CAXI4DMAIIl1I
(
CAXI4DMAIIl1I
)
,
.CAXI4DMAOll1I
(
CAXI4DMAOll1I
)
,
.CAXI4DMAIll1I
(
CAXI4DMAIll1I
)
,
.CAXI4DMAlll1I
(
CAXI4DMAlll1I
)
,
.CAXI4DMAOO01I
(
CAXI4DMAOO01I
)
,
.CAXI4DMAO0l1I
(
CAXI4DMAO0l1I
)
,
.CAXI4DMAl100I
(
CAXI4DMAl100I
)
,
.CAXI4DMAI0l1I
(
CAXI4DMAI0l1I
)
,
.CAXI4DMAl0l1I
(
CAXI4DMAl0l1I
)
,
.CAXI4DMAO1l1I
(
CAXI4DMAO1l1I
)
,
.CAXI4DMAl01Ol
(
CAXI4DMAO011I
)
,
.CAXI4DMAl1OOl
(
CAXI4DMAl1OOl
)
,
.CAXI4DMAl1l1
(
CAXI4DMAl1l1
)
,
.CAXI4DMAO11Ol
(
CAXI4DMAOIOOl
)
,
.CAXI4DMAI11Ol
(
CAXI4DMAIIOOl
)
,
.CAXI4DMAOIOOI
(
CAXI4DMAl111I
)
,
.CAXI4DMAl11Ol
(
CAXI4DMAOOOOl
)
,
.CAXI4DMAOOOIl
(
CAXI4DMAllIOl
)
,
.CAXI4DMAllllI
(
CAXI4DMAO0IOl
)
,
.CAXI4DMAII0OI
(
CAXI4DMAI0IOl
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAlIOOl
)
,
.CAXI4DMAI1IlI
(
CAXI4DMAl0IOl
)
,
.CAXI4DMAIOOIl
(
CAXI4DMAO1IOl
)
,
.CAXI4DMAlOOIl
(
CAXI4DMAI1IOl
)
,
.CAXI4DMAOIOIl
(
CAXI4DMAl1IOl
)
,
.CAXI4DMAIIOIl
(
CAXI4DMAOOlOl
)
,
.CAXI4DMAlIOIl
(
CAXI4DMAIOlOl
)
,
.CAXI4DMAOlOIl
(
CAXI4DMAlOOOl
)
,
.CAXI4DMAIlOIl
(
CAXI4DMAIlIOl
)
)
;
CAXI4DMAllOIl
#
(
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAO1OI
(
CAXI4DMAO1OI
)
,
.NUM_PRI_LVLS
(
NUM_PRI_LVLS
)
,
.CAXI4DMAI1OI
(
CAXI4DMAI1OI
)
,
.PRI_0_NUM_OF_BEATS
(
PRI_0_NUM_OF_BEATS
)
,
.PRI_1_NUM_OF_BEATS
(
PRI_1_NUM_OF_BEATS
)
,
.PRI_2_NUM_OF_BEATS
(
PRI_2_NUM_OF_BEATS
)
,
.PRI_3_NUM_OF_BEATS
(
PRI_3_NUM_OF_BEATS
)
,
.PRI_4_NUM_OF_BEATS
(
PRI_4_NUM_OF_BEATS
)
,
.PRI_5_NUM_OF_BEATS
(
PRI_5_NUM_OF_BEATS
)
,
.PRI_6_NUM_OF_BEATS
(
PRI_6_NUM_OF_BEATS
)
,
.PRI_7_NUM_OF_BEATS
(
PRI_7_NUM_OF_BEATS
)
)
CAXI4DMAO0OIl
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAOOOIl
(
CAXI4DMAllIOl
&
!
CAXI4DMAlI01I
)
,
.CAXI4DMAllllI
(
CAXI4DMAO0IOl
)
,
.CAXI4DMAII0OI
(
CAXI4DMAI0IOl
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAlIOOl
)
,
.CAXI4DMAIOOIl
(
CAXI4DMAO1IOl
)
,
.CAXI4DMAlOOIl
(
CAXI4DMAI1IOl
)
,
.CAXI4DMAOIOIl
(
CAXI4DMAl1IOl
)
,
.CAXI4DMAIIOIl
(
CAXI4DMAOOlOl
)
,
.CAXI4DMAlIOIl
(
CAXI4DMAIOlOl
)
,
.CAXI4DMAI0OIl
(
CAXI4DMAl0IOl
)
,
.CAXI4DMAlII1I
(
CAXI4DMAll00I
)
,
.CAXI4DMAOlI1I
(
CAXI4DMAO000I
)
,
.CAXI4DMAl0OIl
(
CAXI4DMAlO01I
)
,
.CAXI4DMAO1OIl
(
CAXI4DMAII01I
)
,
.CAXI4DMAl011
(
CAXI4DMAl011
)
,
.CAXI4DMAI1OIl
(
CAXI4DMAIIIOl
)
,
.CAXI4DMAl1OIl
(
CAXI4DMAlIIOl
)
,
.CAXI4DMAOlIOl
(
CAXI4DMAOlIOl
)
,
.CAXI4DMAl10Ol
(
CAXI4DMAl10Ol
)
,
.CAXI4DMAO1O1I
(
CAXI4DMAO1O1I
)
,
.CAXI4DMAOIl0I
(
CAXI4DMAIl11I
)
,
.CAXI4DMAOOIIl
(
CAXI4DMAI0OOl
)
,
.CAXI4DMAIllOI
(
CAXI4DMAl0OOl
)
,
.CAXI4DMAO10Ol
(
CAXI4DMAO10Ol
)
,
.CAXI4DMAII
(
CAXI4DMAII
)
,
.CAXI4DMAOl
(
CAXI4DMAOl
)
,
.CAXI4DMAlI
(
CAXI4DMAlI
)
,
.CAXI4DMAll
(
CAXI4DMAll
)
,
.CAXI4DMAO101I
(
CAXI4DMAO101I
)
,
.CAXI4DMAO0
(
CAXI4DMAO0
)
,
.CAXI4DMAlOlOl
(
CAXI4DMAlOlOl
)
,
.CAXI4DMAIIllI
(
CAXI4DMAOIlOl
)
,
.CAXI4DMAO1OOl
(
CAXI4DMAO1OOl
)
)
;
CAXI4DMAIOIIl
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAO1OI
(
CAXI4DMAO1OI
)
,
.AXI4_STREAM_IF
(
AXI4_STREAM_IF
)
)
CAXI4DMAlOIIl
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAIlllI
(
CAXI4DMAIOl1I
)
,
.CAXI4DMAOll0I
(
CAXI4DMAIl01I
)
,
.CAXI4DMAOl0
(
CAXI4DMAOl0
)
,
.CAXI4DMAlI1Ol
(
CAXI4DMAIl0
)
,
.CAXI4DMAl00Ol
(
CAXI4DMAl00Ol
)
,
.CAXI4DMAlOlOl
(
CAXI4DMAlOlOl
)
,
.CAXI4DMAOIlOl
(
CAXI4DMAOIlOl
)
,
.CAXI4DMAOIIIl
(
CAXI4DMAlI0Ol
[
CAXI4DMAl1l1
]
)
,
.CAXI4DMAl01Ol
(
CAXI4DMAO011I
)
,
.CAXI4DMAIIIIl
(
CAXI4DMAIIlOl
)
,
.CAXI4DMAlIIIl
(
CAXI4DMAOllOl
)
,
.CAXI4DMAIOOOl
(
CAXI4DMAIOOOl
)
,
.CAXI4DMAOlOIl
(
CAXI4DMAlOOOl
)
,
.CAXI4DMAOIOOI
(
CAXI4DMAl111I
)
,
.CAXI4DMAl11Ol
(
CAXI4DMAOOOOl
)
,
.CAXI4DMAII0OI
(
CAXI4DMAI0IOl
)
,
.CAXI4DMAIOOIl
(
CAXI4DMAO1IOl
)
,
.CAXI4DMAOOlOl
(
CAXI4DMAOOlOl
)
,
.CAXI4DMAIOlOl
(
CAXI4DMAIOlOl
)
,
.CAXI4DMAOIOOl
(
CAXI4DMAOIOOl
)
,
.CAXI4DMAIIOOl
(
CAXI4DMAIIOOl
)
,
.CAXI4DMAOlIIl
(
CAXI4DMAIlIOl
[
CAXI4DMAOIO1
-
1
:
0
]
)
,
.CAXI4DMAl1l1
(
CAXI4DMAl1l1
)
,
.CAXI4DMAlOllI
(
CAXI4DMAlOllI
)
,
.strDscrptr
(
CAXI4DMAOIllI
)
,
.CAXI4DMAIIllI
(
CAXI4DMAIIllI
)
,
.CAXI4DMAl1IlI
(
CAXI4DMAl1IlI
)
,
.CAXI4DMAOOllI
(
CAXI4DMAOOllI
)
,
.CAXI4DMAIOllI
(
CAXI4DMAIOllI
)
,
.CAXI4DMAl0I0I
(
CAXI4DMAl0I0I
)
,
.intDscrptrNum
(
CAXI4DMAl0l0I
)
)
;
CAXI4DMAIlIIl
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.NUM_PRI_LVLS
(
NUM_PRI_LVLS
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
)
CAXI4DMAllIIl
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAIlllI
(
CAXI4DMAOl0Ol
)
,
.CAXI4DMAO0llI
(
CAXI4DMAO0llI
)
,
.CAXI4DMAI0llI
(
CAXI4DMAI0llI
)
,
.CAXI4DMAlOl1I
(
CAXI4DMAlOl1I
)
,
.CAXI4DMAOIl1I
(
CAXI4DMAOIl1I
)
,
.CAXI4DMAI1l1I
(
CAXI4DMAI1l1I
)
,
.CAXI4DMAIIl1I
(
CAXI4DMAIIl1I
)
,
.CAXI4DMAl1l1I
(
CAXI4DMAl1l1I
)
,
.CAXI4DMAOO01I
(
CAXI4DMAOO01I
)
,
.CAXI4DMAlll1I
(
CAXI4DMAlll1I
)
,
.CAXI4DMAO0l1I
(
CAXI4DMAO0l1I
)
,
.CAXI4DMAl100I
(
CAXI4DMAl100I
)
,
.CAXI4DMAI0l1I
(
CAXI4DMAI0l1I
)
,
.CAXI4DMAl0l1I
(
CAXI4DMAl0l1I
)
,
.CAXI4DMAlIl1I
(
CAXI4DMAlIl1I
)
,
.CAXI4DMAO1l1I
(
CAXI4DMAO1l1I
)
,
.CAXI4DMAI1OOl
(
CAXI4DMAI1OOl
)
,
.CAXI4DMAI1l1
(
CAXI4DMAI1l1
)
,
.CAXI4DMAlOlOl
(
CAXI4DMAlOlOl
)
,
.CAXI4DMAIIllI
(
CAXI4DMAOIlOl
)
,
.CAXI4DMAl1l1
(
CAXI4DMAl1l1
)
,
.CAXI4DMAOOOIl
(
CAXI4DMAIllOl
)
,
.strDscrptr
(
CAXI4DMAO00Ol
)
,
.CAXI4DMAllllI
(
CAXI4DMAI0lOl
)
,
.CAXI4DMAI1IlI
(
CAXI4DMAI00Ol
)
,
.CAXI4DMAIIIIl
(
CAXI4DMAIIlOl
)
,
.CAXI4DMAOIOIl
(
CAXI4DMAlllOl
)
,
.CAXI4DMAlOOIl
(
CAXI4DMAO0lOl
)
,
.CAXI4DMAlIlOl
(
CAXI4DMAlIlOl
)
,
.CAXI4DMAOllOl
(
CAXI4DMAOllOl
)
,
.CAXI4DMAlIOIl
(
CAXI4DMAIOOOl
)
,
.CAXI4DMAO0IIl
(
CAXI4DMAI011I
)
,
.CAXI4DMAI0IIl
(
CAXI4DMAl011I
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAO111I
)
,
.CAXI4DMAII0OI
(
CAXI4DMAI111I
)
,
.CAXI4DMAOIOOI
(
CAXI4DMAl0lOl
)
,
.CAXI4DMAl11Ol
(
CAXI4DMAO1lOl
)
,
.CAXI4DMAOI0Ol
(
CAXI4DMAOI0Ol
)
,
.CAXI4DMAIlOIl
(
CAXI4DMAIl0Ol
)
,
.CAXI4DMAl01Ol
(
CAXI4DMAO011I
)
)
;
CAXI4DMAl0IIl
#
(
.NUM_PRI_LVLS
(
NUM_PRI_LVLS
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAO1OI
(
CAXI4DMAO1OI
)
,
.CAXI4DMAI1OI
(
CAXI4DMAI1OI
)
,
.PRI_0_NUM_OF_BEATS
(
PRI_0_NUM_OF_BEATS
)
,
.PRI_1_NUM_OF_BEATS
(
PRI_1_NUM_OF_BEATS
)
,
.PRI_2_NUM_OF_BEATS
(
PRI_2_NUM_OF_BEATS
)
,
.PRI_3_NUM_OF_BEATS
(
PRI_3_NUM_OF_BEATS
)
,
.PRI_4_NUM_OF_BEATS
(
PRI_4_NUM_OF_BEATS
)
,
.PRI_5_NUM_OF_BEATS
(
PRI_5_NUM_OF_BEATS
)
,
.PRI_6_NUM_OF_BEATS
(
PRI_6_NUM_OF_BEATS
)
,
.PRI_7_NUM_OF_BEATS
(
PRI_7_NUM_OF_BEATS
)
)
CAXI4DMAO1IIl
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAOOOIl
(
CAXI4DMAIllOl
)
,
.CAXI4DMAlIOIl
(
CAXI4DMAIOOOl
)
,
.strDscrptr
(
CAXI4DMAO00Ol
)
,
.CAXI4DMAI1IlI
(
CAXI4DMAI00Ol
)
,
.CAXI4DMAllllI
(
CAXI4DMAI0lOl
)
,
.CAXI4DMAIIIIl
(
CAXI4DMAIIlOl
)
,
.CAXI4DMAOIOIl
(
CAXI4DMAlllOl
)
,
.CAXI4DMAlOOIl
(
CAXI4DMAO0lOl
)
,
.CAXI4DMAI1IIl
(
CAXI4DMAlIlOl
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAO111I
)
,
.CAXI4DMAOO0Ol
(
CAXI4DMAOO0Ol
)
,
.CAXI4DMAl1IIl
(
CAXI4DMAlO0Ol
)
,
.CAXI4DMAOOlIl
(
CAXI4DMAIO01I
)
,
.CAXI4DMAIOlIl
(
CAXI4DMAOI01I
)
,
.CAXI4DMAlOlIl
(
CAXI4DMAlO0
)
,
.CAXI4DMAOIlIl
(
CAXI4DMAOI0
)
,
.CAXI4DMAIIlIl
(
CAXI4DMAll0
)
,
.CAXI4DMAlIlIl
(
CAXI4DMAO00
)
,
.CAXI4DMAOllIl
(
CAXI4DMAOOIOl
)
,
.CAXI4DMAIllIl
(
CAXI4DMAIOIOl
)
,
.CAXI4DMAlllIl
(
CAXI4DMAlOIOl
)
,
.CAXI4DMAO0lIl
(
CAXI4DMAOIIOl
)
,
.CAXI4DMAOO1Ol
(
CAXI4DMAOO1Ol
)
,
.CAXI4DMAI0lIl
(
CAXI4DMAOlOOl
)
,
.CAXI4DMAOllOI
(
CAXI4DMAIlOOl
)
,
.CAXI4DMAl0lIl
(
CAXI4DMAllOOl
)
,
.CAXI4DMAO1lIl
(
CAXI4DMAO0OOl
)
,
.CAXI4DMAI10Ol
(
CAXI4DMAI10Ol
)
,
.CAXI4DMAIOI
(
CAXI4DMAIOI
)
,
.CAXI4DMAOI
(
CAXI4DMAOI
)
,
.CAXI4DMAI0
(
CAXI4DMAI0
)
,
.CAXI4DMAlI0
(
CAXI4DMAOIlOI
)
,
.CAXI4DMAl0
(
CAXI4DMAl0
)
,
.CAXI4DMAI1
(
CAXI4DMAI1
)
,
.CAXI4DMAI101I
(
CAXI4DMAI101I
)
,
.CAXI4DMAll
(
CAXI4DMAOOI
)
,
.CAXI4DMAlOI
(
CAXI4DMAlOI
)
,
.CAXI4DMAOII
(
CAXI4DMAOII
)
,
.CAXI4DMAl00Ol
(
CAXI4DMAl00Ol
)
)
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAII0Ol
<=
2
'b
0
;
end
else
begin
case
(
{
CAXI4DMAl011
,
CAXI4DMAl1lOl
}
)
2
'b
00
:
begin
CAXI4DMAII0Ol
<=
CAXI4DMAII0Ol
;
end
2
'b
01
:
begin
CAXI4DMAII0Ol
[
CAXI4DMAI1l1
]
<=
1
'b
0
;
CAXI4DMAII0Ol
[
!
CAXI4DMAI1l1
]
<=
CAXI4DMAII0Ol
[
!
CAXI4DMAI1l1
]
;
end
2
'b
10
:
begin
CAXI4DMAII0Ol
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAII0Ol
[
!
CAXI4DMAl1l1
]
<=
CAXI4DMAII0Ol
[
!
CAXI4DMAl1l1
]
;
end
2
'b
11
:
begin
if
(
CAXI4DMAI1l1
==
CAXI4DMAl1l1
)
begin
CAXI4DMAII0Ol
<=
CAXI4DMAII0Ol
;
end
else
begin
CAXI4DMAII0Ol
[
CAXI4DMAI1l1
]
<=
1
'b
0
;
CAXI4DMAII0Ol
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
end
end
endcase
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI0Ol
[
0
]
<=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
CAXI4DMAlI0Ol
[
1
]
<=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
end
else
begin
if
(
CAXI4DMAl011
)
begin
CAXI4DMAlI0Ol
[
CAXI4DMAl1l1
]
<=
CAXI4DMAO111
;
end
end
end
assign
CAXI4DMAIO0Ol
=
CAXI4DMAlI0Ol
[
CAXI4DMAl1l1
]
;
assign
CAXI4DMAOO0Ol
=
CAXI4DMAII0Ol
[
CAXI4DMAI1l1
]
;
assign
CAXI4DMAlO0Ol
=
CAXI4DMAlI0Ol
[
CAXI4DMAI1l1
]
;
endmodule
