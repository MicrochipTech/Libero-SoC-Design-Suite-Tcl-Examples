// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAllIOI
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAll1l
,
CAXI4DMAO01l
,
CAXI4DMAI01l
,
CAXI4DMAl01l
,
CAXI4DMAO11l
,
CAXI4DMAI0IOI
,
CAXI4DMAIO01
,
CAXI4DMAlll1
,
CAXI4DMAOOIOI
,
CAXI4DMAOIO0
,
CAXI4DMAIIO0
,
CAXI4DMAO1IOI
,
CAXI4DMAI1IOI
,
CAXI4DMAlI1l
,
CAXI4DMAOIOOI
,
CAXI4DMAl0IOI
)
;
parameter
CAXI4DMAl1OI
=
133
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAO1O1
=
0
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAll1l
;
input
CAXI4DMAO01l
;
input
[
10
:
0
]
CAXI4DMAI01l
;
input
[
31
:
0
]
CAXI4DMAl01l
;
input
[
3
:
0
]
CAXI4DMAO11l
;
input
CAXI4DMAI0IOI
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIO01
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAlll1
;
output
reg
CAXI4DMAOOIOI
;
output
[
31
:
0
]
CAXI4DMAOIO0
;
output
CAXI4DMAIIO0
;
output
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
output
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAI1IOI
;
output
CAXI4DMAlI1l
;
output
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOIOOI
;
output
CAXI4DMAl0IOI
;
localparam
[
4
:
0
]
CAXI4DMAOlIII
=
5
'h
00
;
localparam
[
4
:
0
]
CAXI4DMAIlIII
=
5
'h
04
;
localparam
[
4
:
0
]
CAXI4DMAllIII
=
5
'h
08
;
localparam
[
4
:
0
]
CAXI4DMAO0III
=
5
'h
0C
;
localparam
[
4
:
0
]
CAXI4DMAI0III
=
5
'h
10
;
localparam
[
1
:
0
]
CAXI4DMAOI0l
=
2
'b
01
;
localparam
[
1
:
0
]
CAXI4DMAl0III
=
2
'b
10
;
localparam
[
21
:
0
]
CAXI4DMAlIll
=
22
'b
0000000000000000000001
;
localparam
[
21
:
0
]
CAXI4DMAO1III
=
22
'b
0000000000000000000010
;
localparam
[
21
:
0
]
CAXI4DMAI1III
=
22
'b
0000000000000000000100
;
localparam
[
21
:
0
]
CAXI4DMAl1III
=
22
'b
0000000000000000001000
;
localparam
[
21
:
0
]
CAXI4DMAOOlII
=
22
'b
0000000000000000010000
;
localparam
[
21
:
0
]
CAXI4DMAIOlII
=
22
'b
0000000000000000100000
;
localparam
[
21
:
0
]
CAXI4DMAlOlII
=
22
'b
0000000000000001000000
;
localparam
[
21
:
0
]
CAXI4DMAOIlII
=
22
'b
0000000000000010000000
;
localparam
[
21
:
0
]
CAXI4DMAIIlII
=
22
'b
0000000000000100000000
;
localparam
[
21
:
0
]
CAXI4DMAlIlII
=
22
'b
0000000000001000000000
;
localparam
[
21
:
0
]
CAXI4DMAOllII
=
22
'b
0000000000010000000000
;
localparam
[
21
:
0
]
CAXI4DMAIllII
=
22
'b
0000000000100000000000
;
localparam
[
21
:
0
]
CAXI4DMAlllII
=
22
'b
0000000001000000000000
;
localparam
[
21
:
0
]
CAXI4DMAO0lII
=
22
'b
0000000010000000000000
;
localparam
[
21
:
0
]
CAXI4DMAI0lII
=
22
'b
0000000100000000000000
;
localparam
[
21
:
0
]
CAXI4DMAl0lII
=
22
'b
0000001000000000000000
;
localparam
[
21
:
0
]
CAXI4DMAO1lII
=
22
'b
0000010000000000000000
;
localparam
[
21
:
0
]
CAXI4DMAI1lII
=
22
'b
0000100000000000000000
;
localparam
[
21
:
0
]
CAXI4DMAl1lII
=
22
'b
0001000000000000000000
;
localparam
[
21
:
0
]
CAXI4DMAOO0II
=
22
'b
0010000000000000000000
;
localparam
[
21
:
0
]
CAXI4DMAIO0II
=
22
'b
0100000000000000000000
;
localparam
[
21
:
0
]
CAXI4DMAlO0II
=
22
'b
1000000000000000000000
;
wire
CAXI4DMAOI0II
;
wire
CAXI4DMAII0II
;
wire
CAXI4DMAlI0II
;
wire
CAXI4DMAOl0II
;
wire
CAXI4DMAIl0II
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAll0II
;
reg
[
4
:
0
]
CAXI4DMAOO1
;
reg
[
4
:
0
]
CAXI4DMAO00II
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIO1
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI00II
;
reg
[
31
:
0
]
CAXI4DMAlO1
;
reg
[
31
:
0
]
CAXI4DMAl00II
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAO10II
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAI10II
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAl10II
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOO1II
;
reg
[
1
:
0
]
CAXI4DMAIO1II
;
reg
[
1
:
0
]
CAXI4DMAlO1II
;
wire
[
31
:
0
]
CAXI4DMAOI1II
;
wire
[
31
:
0
]
CAXI4DMAII1II
;
wire
[
31
:
0
]
CAXI4DMAlI1II
;
wire
[
31
:
0
]
CAXI4DMAOl1II
;
wire
[
31
:
0
]
CAXI4DMAIl1II
;
reg
[
21
:
0
]
CAXI4DMAll1II
;
reg
[
21
:
0
]
CAXI4DMAO01II
;
reg
CAXI4DMAI01II
;
reg
CAXI4DMAl01II
;
reg
[
4
:
0
]
CAXI4DMAO11II
;
reg
[
4
:
0
]
CAXI4DMAI11II
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAl11II
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOOOlI
;
reg
[
4
:
0
]
CAXI4DMAIO1l
;
reg
[
4
:
0
]
CAXI4DMAIOOlI
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlI1
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlOOlI
;
reg
CAXI4DMAOIOlI
;
reg
CAXI4DMAIIOlI
;
reg
[
31
:
0
]
CAXI4DMAlIOlI
;
reg
[
31
:
0
]
CAXI4DMAOlOlI
;
reg
CAXI4DMAIIO0
;
reg
CAXI4DMAIlOlI
;
reg
[
31
:
0
]
CAXI4DMAOIO0
;
reg
[
31
:
0
]
CAXI4DMAllOlI
;
reg
CAXI4DMAl0IOI
;
reg
CAXI4DMAO0OlI
;
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAI0OlI
;
wire
CAXI4DMAl0OlI
;
integer
CAXI4DMAO1OlI
;
assign
CAXI4DMAl0OlI
=
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
060
)
&&
(
CAXI4DMAI01l
[
10
:
0
]
<=
11
'h
45C
)
?
CAXI4DMAll1l
:
1
'b
0
;
assign
CAXI4DMAOI0II
=
(
CAXI4DMAI01l
[
4
:
0
]
==
CAXI4DMAOlIII
)
?
CAXI4DMAl0OlI
:
1
'b
0
;
assign
CAXI4DMAII0II
=
(
CAXI4DMAI01l
[
4
:
0
]
==
CAXI4DMAIlIII
)
?
CAXI4DMAl0OlI
:
1
'b
0
;
assign
CAXI4DMAlI0II
=
(
CAXI4DMAI01l
[
4
:
0
]
==
CAXI4DMAllIII
)
?
CAXI4DMAl0OlI
:
1
'b
0
;
assign
CAXI4DMAOl0II
=
(
CAXI4DMAI01l
[
4
:
0
]
==
CAXI4DMAO0III
)
?
CAXI4DMAl0OlI
:
1
'b
0
;
assign
CAXI4DMAIl0II
=
(
CAXI4DMAI01l
[
4
:
0
]
==
CAXI4DMAI0III
)
?
CAXI4DMAl0OlI
:
1
'b
0
;
assign
CAXI4DMAll0II
=
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
8
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
9
)
)
?
5
'd
1
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
A
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
B
)
)
?
5
'd
2
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
C
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
D
)
)
?
5
'd
3
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
E
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
F
)
)
?
5
'd
4
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
10
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
11
)
)
?
5
'd
5
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
12
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
13
)
)
?
5
'd
6
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
14
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
15
)
)
?
5
'd
7
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
16
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
17
)
)
?
5
'd
8
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
18
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
19
)
)
?
5
'd
9
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
1A
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
1B
)
)
?
5
'd
10
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
1C
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
1D
)
)
?
5
'd
11
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
1E
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
1F
)
)
?
5
'd
12
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
20
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
21
)
)
?
5
'd
13
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
22
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
23
)
)
?
5
'd
14
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
24
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
25
)
)
?
5
'd
15
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
26
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
27
)
)
?
5
'd
16
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
28
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
29
)
)
?
5
'd
17
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
2A
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
2B
)
)
?
5
'd
18
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
2C
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
2D
)
)
?
5
'd
19
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
2E
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
2F
)
)
?
5
'd
20
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
30
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
31
)
)
?
5
'd
21
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
32
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
33
)
)
?
5
'd
22
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
34
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
35
)
)
?
5
'd
23
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
36
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
37
)
)
?
5
'd
24
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
38
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
39
)
)
?
5
'd
25
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
3A
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
3B
)
)
?
5
'd
26
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
3C
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
3D
)
)
?
5
'd
27
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
3E
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
3F
)
)
?
5
'd
28
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
40
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
41
)
)
?
5
'd
29
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
42
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
43
)
)
?
5
'd
30
:
(
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
44
)
||
(
CAXI4DMAI01l
[
10
:
4
]
==
7
'h
45
)
)
?
5
'd
31
:
5
'd
0
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOO1
<=
5
'b
0
;
end
else
begin
CAXI4DMAOO1
<=
CAXI4DMAO00II
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO1
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIO1
<=
CAXI4DMAI00II
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlO1
<=
32
'd
0
;
end
else
begin
CAXI4DMAlO1
<=
CAXI4DMAl00II
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI1
<=
32
'd
0
;
end
else
begin
CAXI4DMAlI1
<=
CAXI4DMAlOOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO1l
<=
5
'd
0
;
end
else
begin
CAXI4DMAIO1l
<=
CAXI4DMAIOOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI01II
<=
1
'b
0
;
end
else
begin
CAXI4DMAI01II
<=
CAXI4DMAl01II
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO11II
<=
5
'b
0
;
end
else
begin
CAXI4DMAO11II
<=
CAXI4DMAI11II
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl11II
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAl11II
<=
CAXI4DMAOOOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIOlI
<=
1
'b
0
;
end
else
begin
CAXI4DMAOIOlI
<=
CAXI4DMAIIOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlIOlI
<=
32
'b
0
;
end
else
begin
CAXI4DMAlIOlI
<=
CAXI4DMAOlOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIIO0
<=
1
'b
0
;
end
else
begin
CAXI4DMAIIO0
<=
CAXI4DMAIlOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIO0
<=
32
'b
0
;
end
else
begin
CAXI4DMAOIO0
<=
CAXI4DMAllOlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0IOI
<=
1
'b
0
;
end
else
begin
CAXI4DMAl0IOI
<=
CAXI4DMAO0OlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO1IOI
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAO1IOI
<=
CAXI4DMAI0OlI
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO1II
<=
CAXI4DMAOI0l
;
end
else
begin
CAXI4DMAIO1II
<=
CAXI4DMAlO1II
;
end
end
always
@
(
*
)
begin
CAXI4DMAO00II
<=
5
'b
0
;
CAXI4DMAI00II
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAl00II
<=
32
'b
0
;
CAXI4DMAOOIOI
<=
1
'b
0
;
CAXI4DMAl01II
<=
1
'b
0
;
CAXI4DMAI11II
<=
5
'b
0
;
CAXI4DMAOOOlI
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
case
(
CAXI4DMAIO1II
)
CAXI4DMAOI0l
:
begin
if
(
(
CAXI4DMAOI0II
|
CAXI4DMAII0II
|
CAXI4DMAlI0II
|
CAXI4DMAOl0II
|
CAXI4DMAIl0II
)
&&
CAXI4DMAO01l
)
begin
if
(
CAXI4DMAO11l
!=
4
'h
F
)
begin
CAXI4DMAl01II
<=
1
'b
1
;
CAXI4DMAI11II
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAOOOlI
<=
CAXI4DMAll0II
;
CAXI4DMAlO1II
<=
CAXI4DMAl0III
;
end
else
begin
CAXI4DMAO00II
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAI00II
<=
CAXI4DMAll0II
;
CAXI4DMAl00II
<=
CAXI4DMAl01l
;
CAXI4DMAOOIOI
<=
1
'b
1
;
CAXI4DMAlO1II
<=
CAXI4DMAOI0l
;
end
end
else
begin
CAXI4DMAlO1II
<=
CAXI4DMAOI0l
;
end
end
CAXI4DMAl0III
:
begin
if
(
CAXI4DMAOIOlI
)
begin
CAXI4DMAO00II
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAI00II
<=
CAXI4DMAll0II
;
CAXI4DMAl00II
[
31
:
24
]
<=
(
CAXI4DMAO11l
[
3
]
)
?
CAXI4DMAl01l
[
31
:
24
]
:
CAXI4DMAlIOlI
[
31
:
24
]
;
CAXI4DMAl00II
[
23
:
16
]
<=
(
CAXI4DMAO11l
[
2
]
)
?
CAXI4DMAl01l
[
23
:
16
]
:
CAXI4DMAlIOlI
[
23
:
16
]
;
CAXI4DMAl00II
[
15
:
8
]
<=
(
CAXI4DMAO11l
[
1
]
)
?
CAXI4DMAl01l
[
15
:
8
]
:
CAXI4DMAlIOlI
[
15
:
8
]
;
CAXI4DMAl00II
[
7
:
0
]
<=
(
CAXI4DMAO11l
[
0
]
)
?
CAXI4DMAl01l
[
7
:
0
]
:
CAXI4DMAlIOlI
[
7
:
0
]
;
CAXI4DMAOOIOI
<=
1
'b
1
;
CAXI4DMAlO1II
<=
CAXI4DMAOI0l
;
end
else
begin
CAXI4DMAl01II
<=
1
'b
1
;
CAXI4DMAI11II
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAOOOlI
<=
CAXI4DMAll0II
;
CAXI4DMAlO1II
<=
CAXI4DMAl0III
;
end
end
default
:
begin
CAXI4DMAlO1II
<=
CAXI4DMAOI0l
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO10II
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
end
else
begin
if
(
CAXI4DMAOI0II
&
CAXI4DMAO11l
[
1
]
&
CAXI4DMAl01l
[
15
]
&
CAXI4DMAOOIOI
)
begin
CAXI4DMAO10II
[
CAXI4DMAll0II
]
<=
1
'b
1
;
end
else
if
(
CAXI4DMAOOIOI
&&
(
(
(
CAXI4DMAIl0II
|
CAXI4DMAOl0II
|
CAXI4DMAlI0II
|
CAXI4DMAII0II
)
&
~
CAXI4DMAOI0II
)
||
(
CAXI4DMAOI0II
&
(
~
CAXI4DMAO11l
[
1
]
|
(
CAXI4DMAO11l
[
1
]
&
~
CAXI4DMAl01l
[
15
]
)
)
)
)
)
begin
CAXI4DMAO10II
[
CAXI4DMAll0II
]
<=
1
'b
0
;
end
end
end
assign
CAXI4DMAlI1l
=
CAXI4DMAO10II
[
CAXI4DMAIO01
]
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
for
(
CAXI4DMAO1OlI
=
0
;
CAXI4DMAO1OlI
<
NUM_INT_BDS
;
CAXI4DMAO1OlI
=
CAXI4DMAO1OlI
+
1
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI10II
[
CAXI4DMAO1OlI
]
<=
1
'b
0
;
end
else
begin
if
(
CAXI4DMAOI0II
&
CAXI4DMAO11l
[
1
]
&
CAXI4DMAOOIOI
&
(
CAXI4DMAll0II
==
CAXI4DMAO1OlI
)
)
begin
CAXI4DMAI10II
[
CAXI4DMAO1OlI
]
<=
CAXI4DMAl01l
[
13
]
;
end
else
begin
CAXI4DMAI10II
[
CAXI4DMAO1OlI
]
<=
CAXI4DMAI10II
[
CAXI4DMAO1OlI
]
&
~
CAXI4DMAlll1
[
CAXI4DMAO1OlI
]
;
end
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
for
(
CAXI4DMAO1OlI
=
0
;
CAXI4DMAO1OlI
<
NUM_INT_BDS
;
CAXI4DMAO1OlI
=
CAXI4DMAO1OlI
+
1
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10II
[
CAXI4DMAO1OlI
]
<=
1
'b
0
;
end
else
begin
if
(
CAXI4DMAOI0II
&
CAXI4DMAO11l
[
1
]
&
CAXI4DMAOOIOI
&
(
CAXI4DMAll0II
==
CAXI4DMAO1OlI
)
)
begin
CAXI4DMAl10II
[
CAXI4DMAO1OlI
]
<=
CAXI4DMAl01l
[
14
]
;
end
else
begin
CAXI4DMAl10II
[
CAXI4DMAO1OlI
]
<=
CAXI4DMAl10II
[
CAXI4DMAO1OlI
]
&
~
CAXI4DMAlll1
[
CAXI4DMAO1OlI
]
;
end
end
end
end
assign
CAXI4DMAI1IOI
=
CAXI4DMAI10II
&
CAXI4DMAl10II
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOO1II
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
end
else
begin
if
(
CAXI4DMAOI0II
&
CAXI4DMAO11l
[
1
]
&
CAXI4DMAOOIOI
)
begin
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
<=
CAXI4DMAl01l
[
10
]
;
end
else
begin
CAXI4DMAOO1II
<=
CAXI4DMAOO1II
;
end
end
end
assign
CAXI4DMAOIOOI
=
CAXI4DMAOO1II
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAll1II
<=
CAXI4DMAlIll
;
end
else
begin
CAXI4DMAll1II
<=
CAXI4DMAO01II
;
end
end
always
@
(
*
)
begin
CAXI4DMAIOOlI
<=
{
5
{
1
'b
0
}
}
;
CAXI4DMAlOOlI
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAIIOlI
<=
1
'b
0
;
CAXI4DMAOlOlI
<=
32
'b
0
;
CAXI4DMAIlOlI
<=
1
'b
0
;
CAXI4DMAllOlI
<=
32
'b
0
;
CAXI4DMAO0OlI
<=
1
'b
0
;
CAXI4DMAI0OlI
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
case
(
CAXI4DMAll1II
)
CAXI4DMAlIll
:
begin
if
(
CAXI4DMAI01II
)
begin
CAXI4DMAIOOlI
<=
CAXI4DMAO11II
;
CAXI4DMAlOOlI
<=
CAXI4DMAl11II
;
CAXI4DMAO01II
<=
CAXI4DMAO1III
;
end
else
if
(
(
CAXI4DMAIl0II
|
CAXI4DMAOl0II
|
CAXI4DMAlI0II
|
CAXI4DMAII0II
|
CAXI4DMAOI0II
)
&&
~
CAXI4DMAO01l
)
begin
CAXI4DMAIOOlI
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAlOOlI
<=
CAXI4DMAll0II
;
CAXI4DMAO01II
<=
CAXI4DMAO1lII
;
end
else
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAOIlII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAlIll
;
end
end
CAXI4DMAO1III
:
begin
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAl1III
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAI1III
;
end
end
CAXI4DMAI1III
:
begin
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAIOlII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAOOlII
;
end
end
CAXI4DMAl1III
:
begin
CAXI4DMAO01II
<=
CAXI4DMAlOlII
;
end
CAXI4DMAOOlII
:
begin
CAXI4DMAIIOlI
<=
1
'b
1
;
if
(
CAXI4DMAO11II
[
0
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAOI1II
;
end
else
if
(
CAXI4DMAO11II
[
1
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAII1II
;
end
else
if
(
CAXI4DMAO11II
[
2
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAlI1II
;
end
else
if
(
CAXI4DMAO11II
[
3
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAOl1II
;
end
else
if
(
CAXI4DMAO11II
[
4
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAIl1II
;
end
else
begin
CAXI4DMAOlOlI
<=
32
'b
0
;
end
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAOIlII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAlIll
;
end
end
CAXI4DMAIOlII
:
begin
CAXI4DMAIIOlI
<=
1
'b
1
;
if
(
CAXI4DMAO11II
[
0
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAOI1II
;
end
else
if
(
CAXI4DMAO11II
[
1
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAII1II
;
end
else
if
(
CAXI4DMAO11II
[
2
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAlI1II
;
end
else
if
(
CAXI4DMAO11II
[
3
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAOl1II
;
end
else
if
(
CAXI4DMAO11II
[
4
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAIl1II
;
end
else
begin
CAXI4DMAOlOlI
<=
32
'b
0
;
end
CAXI4DMAO01II
<=
CAXI4DMAIIlII
;
end
CAXI4DMAlOlII
:
begin
CAXI4DMAIIOlI
<=
1
'b
1
;
if
(
CAXI4DMAO11II
[
0
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAOI1II
;
end
else
if
(
CAXI4DMAO11II
[
1
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAII1II
;
end
else
if
(
CAXI4DMAO11II
[
2
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAlI1II
;
end
else
if
(
CAXI4DMAO11II
[
3
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAOl1II
;
end
else
if
(
CAXI4DMAO11II
[
4
]
)
begin
CAXI4DMAOlOlI
<=
CAXI4DMAIl1II
;
end
else
begin
CAXI4DMAOlOlI
<=
32
'b
0
;
end
CAXI4DMAO01II
<=
CAXI4DMAIllII
;
end
CAXI4DMAOIlII
:
begin
if
(
CAXI4DMAI01II
)
begin
CAXI4DMAIOOlI
<=
CAXI4DMAO11II
;
CAXI4DMAlOOlI
<=
CAXI4DMAl11II
;
CAXI4DMAO01II
<=
CAXI4DMAlIlII
;
end
else
if
(
(
CAXI4DMAIl0II
|
CAXI4DMAOl0II
|
CAXI4DMAlI0II
|
CAXI4DMAII0II
|
CAXI4DMAOI0II
)
&&
~
CAXI4DMAO01l
)
begin
CAXI4DMAIOOlI
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAlOOlI
<=
CAXI4DMAll0II
;
CAXI4DMAO01II
<=
CAXI4DMAOllII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAIIlII
;
end
end
CAXI4DMAIIlII
:
begin
if
(
CAXI4DMAI01II
)
begin
CAXI4DMAIOOlI
<=
CAXI4DMAO11II
;
CAXI4DMAlOOlI
<=
CAXI4DMAl11II
;
CAXI4DMAO01II
<=
CAXI4DMAlllII
;
end
else
if
(
(
CAXI4DMAIl0II
|
CAXI4DMAOl0II
|
CAXI4DMAlI0II
|
CAXI4DMAII0II
|
CAXI4DMAOI0II
)
&&
~
CAXI4DMAO01l
)
begin
CAXI4DMAIOOlI
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAlOOlI
<=
CAXI4DMAll0II
;
CAXI4DMAO01II
<=
CAXI4DMAI0lII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAIllII
;
end
end
CAXI4DMAlIlII
:
begin
CAXI4DMAO01II
<=
CAXI4DMAO0lII
;
end
CAXI4DMAOllII
:
begin
CAXI4DMAO01II
<=
CAXI4DMAl0lII
;
end
CAXI4DMAIllII
:
begin
CAXI4DMAO0OlI
<=
1
'b
1
;
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
if
(
CAXI4DMAI01II
)
begin
CAXI4DMAIOOlI
<=
CAXI4DMAO11II
;
CAXI4DMAlOOlI
<=
CAXI4DMAl11II
;
CAXI4DMAO01II
<=
CAXI4DMAO1III
;
end
else
if
(
(
CAXI4DMAIl0II
|
CAXI4DMAOl0II
|
CAXI4DMAlI0II
|
CAXI4DMAII0II
|
CAXI4DMAOI0II
)
&&
~
CAXI4DMAO01l
)
begin
CAXI4DMAIOOlI
<=
{
CAXI4DMAIl0II
,
CAXI4DMAOl0II
,
CAXI4DMAlI0II
,
CAXI4DMAII0II
,
CAXI4DMAOI0II
}
;
CAXI4DMAlOOlI
<=
CAXI4DMAll0II
;
CAXI4DMAO01II
<=
CAXI4DMAO1lII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAlIll
;
end
end
CAXI4DMAlllII
:
begin
CAXI4DMAO0OlI
<=
1
'b
1
;
CAXI4DMAO01II
<=
CAXI4DMAI1III
;
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
CAXI4DMAO0lII
:
begin
CAXI4DMAO0OlI
<=
1
'b
1
;
CAXI4DMAO01II
<=
CAXI4DMAOOlII
;
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
CAXI4DMAI0lII
:
begin
CAXI4DMAO0OlI
<=
1
'b
1
;
CAXI4DMAO01II
<=
CAXI4DMAI1lII
;
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
CAXI4DMAl0lII
:
begin
CAXI4DMAO0OlI
<=
1
'b
1
;
CAXI4DMAO01II
<=
CAXI4DMAOO0II
;
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAI0OlI
<=
{
CAXI4DMAIl1II
,
CAXI4DMAOl1II
,
CAXI4DMAlI1II
,
CAXI4DMAII1II
[
23
:
0
]
,
CAXI4DMAI1IOI
[
CAXI4DMAIO01
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAIO01
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
CAXI4DMAO1lII
:
begin
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAl1lII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAI1lII
;
end
end
CAXI4DMAI1lII
:
begin
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAIO0II
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAOO0II
;
end
end
CAXI4DMAl1lII
:
begin
CAXI4DMAO01II
<=
CAXI4DMAlO0II
;
end
CAXI4DMAOO0II
:
begin
CAXI4DMAIlOlI
<=
1
'b
1
;
if
(
CAXI4DMAOI0II
)
begin
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAllOlI
<=
{
CAXI4DMAOI1II
[
31
:
16
]
,
CAXI4DMAO10II
[
CAXI4DMAll0II
]
,
CAXI4DMAl10II
[
CAXI4DMAll0II
]
,
CAXI4DMAI10II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAllOlI
<=
{
CAXI4DMAOI1II
[
31
:
16
]
,
CAXI4DMAO10II
[
CAXI4DMAll0II
]
,
CAXI4DMAl10II
[
CAXI4DMAll0II
]
,
CAXI4DMAI10II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
else
if
(
CAXI4DMAII0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAII1II
;
end
else
if
(
CAXI4DMAlI0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAlI1II
;
end
else
if
(
CAXI4DMAOl0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAOl1II
;
end
else
if
(
CAXI4DMAIl0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAIl1II
;
end
else
begin
CAXI4DMAllOlI
<=
32
'b
0
;
end
if
(
CAXI4DMAI0IOI
)
begin
CAXI4DMAIOOlI
<=
5
'b
11111
;
CAXI4DMAlOOlI
<=
CAXI4DMAIO01
;
CAXI4DMAO01II
<=
CAXI4DMAOIlII
;
end
else
begin
CAXI4DMAO01II
<=
CAXI4DMAlIll
;
end
end
CAXI4DMAIO0II
:
begin
CAXI4DMAIlOlI
<=
1
'b
1
;
if
(
CAXI4DMAOI0II
)
begin
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAllOlI
<=
{
CAXI4DMAOI1II
[
31
:
16
]
,
CAXI4DMAO10II
[
CAXI4DMAll0II
]
,
CAXI4DMAl10II
[
CAXI4DMAll0II
]
,
CAXI4DMAI10II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAllOlI
<=
{
CAXI4DMAOI1II
[
31
:
16
]
,
CAXI4DMAO10II
[
CAXI4DMAll0II
]
,
CAXI4DMAl10II
[
CAXI4DMAll0II
]
,
CAXI4DMAI10II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
else
if
(
CAXI4DMAII0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAII1II
;
end
else
if
(
CAXI4DMAlI0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAlI1II
;
end
else
if
(
CAXI4DMAOl0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAOl1II
;
end
else
if
(
CAXI4DMAIl0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAIl1II
;
end
else
begin
CAXI4DMAllOlI
<=
32
'b
0
;
end
CAXI4DMAO01II
<=
CAXI4DMAIIlII
;
end
CAXI4DMAlO0II
:
begin
CAXI4DMAIlOlI
<=
1
'b
1
;
if
(
CAXI4DMAOI0II
)
begin
if
(
CAXI4DMAO1O1
==
1
)
begin
CAXI4DMAllOlI
<=
{
CAXI4DMAOI1II
[
31
:
16
]
,
CAXI4DMAO10II
[
CAXI4DMAll0II
]
,
CAXI4DMAl10II
[
CAXI4DMAll0II
]
,
CAXI4DMAI10II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
9
:
0
]
}
;
end
else
begin
CAXI4DMAllOlI
<=
{
CAXI4DMAOI1II
[
31
:
16
]
,
CAXI4DMAO10II
[
CAXI4DMAll0II
]
,
CAXI4DMAl10II
[
CAXI4DMAll0II
]
,
CAXI4DMAI10II
[
CAXI4DMAll0II
]
,
CAXI4DMAOI1II
[
12
:
11
]
,
CAXI4DMAOO1II
[
CAXI4DMAll0II
]
,
{
6
{
1
'b
0
}
}
,
CAXI4DMAOI1II
[
3
:
0
]
}
;
end
end
else
if
(
CAXI4DMAII0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAII1II
;
end
else
if
(
CAXI4DMAlI0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAlI1II
;
end
else
if
(
CAXI4DMAOl0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAOl1II
;
end
else
if
(
CAXI4DMAIl0II
)
begin
CAXI4DMAllOlI
<=
CAXI4DMAIl1II
;
end
else
begin
CAXI4DMAllOlI
<=
32
'b
0
;
end
CAXI4DMAO01II
<=
CAXI4DMAIllII
;
end
default
:
begin
CAXI4DMAO01II
<=
CAXI4DMAlIll
;
end
endcase
end
CAXI4DMAI1OlI
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl1OlI
(
1
'b
1
)
)
CAXI4DMAOOIlI
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAOO1
(
CAXI4DMAOO1
[
0
]
)
,
.CAXI4DMAIO1
(
CAXI4DMAIO1
)
,
.CAXI4DMAlO1
(
CAXI4DMAlO1
)
,
.CAXI4DMAIO1l
(
CAXI4DMAIO1l
[
0
]
)
,
.CAXI4DMAlI1
(
CAXI4DMAlI1
)
,
.CAXI4DMAI1Il
(
CAXI4DMAOI1II
)
)
;
CAXI4DMAI1OlI
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl1OlI
(
1
'b
1
)
)
CAXI4DMAIOIlI
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAOO1
(
CAXI4DMAOO1
[
1
]
)
,
.CAXI4DMAIO1
(
CAXI4DMAIO1
)
,
.CAXI4DMAlO1
(
CAXI4DMAlO1
)
,
.CAXI4DMAIO1l
(
CAXI4DMAIO1l
[
1
]
)
,
.CAXI4DMAlI1
(
CAXI4DMAlI1
)
,
.CAXI4DMAI1Il
(
CAXI4DMAII1II
)
)
;
CAXI4DMAI1OlI
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl1OlI
(
1
'b
1
)
)
CAXI4DMAlOIlI
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAOO1
(
CAXI4DMAOO1
[
2
]
)
,
.CAXI4DMAIO1
(
CAXI4DMAIO1
)
,
.CAXI4DMAlO1
(
CAXI4DMAlO1
)
,
.CAXI4DMAIO1l
(
CAXI4DMAIO1l
[
2
]
)
,
.CAXI4DMAlI1
(
CAXI4DMAlI1
)
,
.CAXI4DMAI1Il
(
CAXI4DMAlI1II
)
)
;
CAXI4DMAI1OlI
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl1OlI
(
1
'b
1
)
)
CAXI4DMAOIIlI
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAOO1
(
CAXI4DMAOO1
[
3
]
)
,
.CAXI4DMAIO1
(
CAXI4DMAIO1
)
,
.CAXI4DMAlO1
(
CAXI4DMAlO1
)
,
.CAXI4DMAIO1l
(
CAXI4DMAIO1l
[
3
]
)
,
.CAXI4DMAlI1
(
CAXI4DMAlI1
)
,
.CAXI4DMAI1Il
(
CAXI4DMAOl1II
)
)
;
CAXI4DMAI1OlI
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl1OlI
(
1
'b
1
)
)
CAXI4DMAIIIlI
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAOO1
(
CAXI4DMAOO1
[
4
]
)
,
.CAXI4DMAIO1
(
CAXI4DMAIO1
)
,
.CAXI4DMAlO1
(
CAXI4DMAlO1
)
,
.CAXI4DMAIO1l
(
CAXI4DMAIO1l
[
4
]
)
,
.CAXI4DMAlI1
(
CAXI4DMAlI1
)
,
.CAXI4DMAI1Il
(
CAXI4DMAIl1II
)
)
;
endmodule
