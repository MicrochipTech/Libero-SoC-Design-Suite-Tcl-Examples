`timescale 1 ns/100 ps
// Version: v12.6 12.900.20.6


module ACT_UNIQUE_prbsgen_parallel_fab(
       prbsgen_parallel_fab_0_prbs_out_msb_o_0,
       current_state_0,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G
    );
output [7:0] prbsgen_parallel_fab_0_prbs_out_msb_o_0;
input  current_state_0;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;

    wire [7:0] s_prbsin_Z;
    wire GND, VCC;
    
    GND GND_Z (.Y(GND));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[1]  (.A(s_prbsin_Z[7]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7]), .Y(s_prbsin_Z[1]));
    VCC VCC_Z (.Y(VCC));
    SLE \prbs_out_o[2]  (.D(s_prbsin_Z[2]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5]));
    SLE \prbs_out_o[1]  (.D(s_prbsin_Z[1]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[5]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4]), .Y(s_prbsin_Z[5]));
    SLE \prbs_out_o[7]  (.D(s_prbsin_Z[7]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[0]));
    SLE \prbs_out_o[6]  (.D(s_prbsin_Z[6]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[7]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2]), .Y(s_prbsin_Z[7]));
    SLE \prbs_out_o[5]  (.D(s_prbsin_Z[5]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[0]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3]), .Y(s_prbsin_Z[0]));
    SLE \prbs_out_o[4]  (.D(s_prbsin_Z[4]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3]));
    SLE \prbs_out_o[0]  (.D(s_prbsin_Z[0]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[2]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7]), .Y(s_prbsin_Z[2]));
    SLE \prbs_out_o[3]  (.D(s_prbsin_Z[3]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(current_state_0), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[4]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5]), .Y(s_prbsin_Z[4]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[6]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3]), .Y(s_prbsin_Z[6]));
    CFG2 #( .INIT(4'h6) )  \s_prbsin[3]  (.A(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5]), .B(
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6]), .Y(s_prbsin_Z[3]));
    
endmodule


module PLL_BCLKSCLKALIGN_Z5(
       current_state_RNI00O7_Y_0,
       current_state_0,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX,
       N_386_i,
       PLL_LOCK_0,
       COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL,
       N_81,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       DB_OUT
    );
output current_state_RNI00O7_Y_0;
output current_state_0;
input  [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
output N_386_i;
input  PLL_LOCK_0;
output COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL;
output N_81;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;
input  DB_OUT;

    wire [4:0] dly_cnt_Z;
    wire [3:0] reset_cycle_count_Z;
    wire [2:2] rotate_count_Z;
    wire [2:2] rotate_count_4;
    wire [3:0] bclk_igear_rx_reg_Z;
    wire [15:0] current_state_Z;
    wire [15:0] current_state_ns;
    wire [9:0] transition_check_counter_Z;
    wire [8:0] transition_check_counter_s;
    wire [9:9] transition_check_counter_s_Z;
    wire [6:0] vcophsel_bclk_Z;
    wire [6:0] vcophsel_bclk_s;
    wire [0:0] transition_check_counter_cry_cy_S;
    wire [0:0] transition_check_counter_cry_cy_Y;
    wire [8:0] transition_check_counter_cry_Z;
    wire [8:0] transition_check_counter_cry_Y;
    wire [9:9] transition_check_counter_s_FCO;
    wire [9:9] transition_check_counter_s_Y;
    wire [1:1] current_state_RNI00O7_S;
    wire [5:0] vcophsel_bclk_cry;
    wire [0:0] vcophsel_bclk_RNIRNHR_Y;
    wire [1:1] vcophsel_bclk_RNINGBF1_Y;
    wire [2:2] vcophsel_bclk_RNIKA532_Y;
    wire [3:3] vcophsel_bclk_RNII5VM2_Y;
    wire [4:4] vcophsel_bclk_RNIH1PA3_Y;
    wire [6:6] vcophsel_bclk_RNO_FCO;
    wire [6:6] vcophsel_bclk_RNO_Y;
    wire [5:5] vcophsel_bclk_RNIHUIU3_Y;
    wire [0:0] current_state_ns_a2_0_a2_5_Z;
    wire [0:0] current_state_ns_a2_0_a2_3_Z;
    wire [4:4] current_state_ns_a2_1_6_Z;
    wire [4:4] current_state_ns_a2_1_5_Z;
    wire [0:0] current_state_ns_a2_0_a2_7_Z;
    wire VCC, N_23, N_97_i, GND, N_88_i, N_91_i, N_82_i, N_85_i, 
        N_47_i, next_state43_0, N_77_i, next_state43_1, N_78_i_i, 
        N_374_i, N_53_i, N_51_i, N_49_i, N_315_i_0, N_59_i, N_64, 
        N_38_i, N_281_i, N_41_i, N_284_i, N_287_i, N_354_i, 
        transition_detected_Z, transition_detected_3, N_126_i, 
        transition_check_counter_cry_cy, vcophsel_bclk_cry_cy, N_69, 
        N_62_i, N_144, un4_transition_detected_1, 
        un4_transition_detected_0, un1_vcophsel_bclk_1_4_Z, N_145, 
        un8_transition_detected, un10_transition_detected, N_68, N_72, 
        un1_vcophsel_bclk_1_Z, N_212, un1_rst_clk_align_trng_1_0_0_Z, 
        N_76, N_436, N_435, N_434, N_412, N_411, N_410, N_409, N_408, 
        N_407, N_406, N_405, N_404, N_403, N_402, N_401, N_400, N_399, 
        N_398, N_397, N_396, N_395, N_394, N_393, N_46, N_45, N_44, 
        N_43, N_42, N_41, N_40, N_39, N_38, N_37, N_36, N_35, N_34, 
        N_33, N_32, N_31, N_30, N_29, N_28, N_27, N_26, N_25, N_24, 
        N_23_0, N_22, N_21, N_20, N_19, N_18, N_17, N_16, N_15, N_7;
    
    SLE \rotate_count[0]  (.D(N_77_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(next_state43_0));
    CFG3 #( .INIT(8'h01) )  \current_state_ns_a2_0_a2_3[0]  (.A(
        current_state_Z[15]), .B(PLL_LOCK_0), .C(current_state_Z[3]), 
        .Y(current_state_ns_a2_0_a2_3_Z[0]));
    CFG4 #( .INIT(16'h0C06) )  \reset_cycle_count_RNO[3]  (.A(
        reset_cycle_count_Z[2]), .B(reset_cycle_count_Z[3]), .C(
        un1_rst_clk_align_trng_1_0_0_Z), .D(N_72), .Y(N_47_i));
    SLE \transition_check_counter[2]  (.D(
        transition_check_counter_s[2]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[2]));
    SLE \transition_check_counter[7]  (.D(
        transition_check_counter_s[7]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[7]));
    SLE \dly_cnt[2]  (.D(N_23), .CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(
        N_97_i), .ALn(DB_OUT), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(dly_cnt_Z[2]));
    CFG4 #( .INIT(16'hFFFE) )  \dly_cnt_RNIARNS[3]  (.A(dly_cnt_Z[3]), 
        .B(dly_cnt_Z[2]), .C(dly_cnt_Z[1]), .D(dly_cnt_Z[0]), .Y(N_69));
    ARI1 #( .INIT(20'h45500) )  \transition_check_counter_cry_cy[0]  (
        .A(VCC), .B(current_state_Z[5]), .C(GND), .D(GND), .FCI(VCC), 
        .S(transition_check_counter_cry_cy_S[0]), .Y(
        transition_check_counter_cry_cy_Y[0]), .FCO(
        transition_check_counter_cry_cy));
    CFG4 #( .INIT(16'h1000) )  \current_state_ns_a2_0_a2[9]  (.A(
        next_state43_1), .B(next_state43_0), .C(rotate_count_Z[2]), .D(
        current_state_Z[6]), .Y(current_state_ns[9]));
    SLE \current_state[3]  (.D(current_state_Z[2]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_315_i_0), .ALn(DB_OUT), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        current_state_Z[3]));
    SLE \vcophsel_bclk[2]  (.D(vcophsel_bclk_s[2]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[2]));
    CFG3 #( .INIT(8'h41) )  \reset_cycle_count_RNO[2]  (.A(
        un1_rst_clk_align_trng_1_0_0_Z), .B(reset_cycle_count_Z[2]), 
        .C(N_72), .Y(N_49_i));
    SLE \vcophsel_bclk[0]  (.D(vcophsel_bclk_s[0]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[0]));
    CFG2 #( .INIT(4'h6) )  \rotate_count_RNO[0]  (.A(
        current_state_Z[8]), .B(next_state43_0), .Y(N_77_i));
    CFG4 #( .INIT(16'h0001) )  \current_state_ns_a2_1_5[4]  (.A(
        transition_check_counter_Z[9]), .B(
        transition_check_counter_Z[8]), .C(
        transition_check_counter_Z[5]), .D(
        transition_check_counter_Z[4]), .Y(
        current_state_ns_a2_1_5_Z[4]));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNIRNHR[0]  (.A(VCC), 
        .B(current_state_Z[1]), .C(vcophsel_bclk_Z[0]), .D(GND), .FCI(
        vcophsel_bclk_cry_cy), .S(vcophsel_bclk_s[0]), .Y(
        vcophsel_bclk_RNIRNHR_Y[0]), .FCO(vcophsel_bclk_cry[0]));
    CFG4 #( .INIT(16'hC0D5) )  \current_state_ns_0[5]  (.A(N_212), .B(
        current_state_Z[3]), .C(N_315_i_0), .D(N_76), .Y(
        current_state_ns[5]));
    SLE \transition_check_counter[0]  (.D(
        transition_check_counter_s[0]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[0]));
    CFG4 #( .INIT(16'hFFFE) )  \register_rx.un10_transition_detected  
        (.A(bclk_igear_rx_reg_Z[3]), .B(bclk_igear_rx_reg_Z[2]), .C(
        bclk_igear_rx_reg_Z[1]), .D(bclk_igear_rx_reg_Z[0]), .Y(
        un10_transition_detected));
    SLE \rotate_count[2]  (.D(rotate_count_4[2]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(rotate_count_Z[2]));
    SLE \dly_cnt[0]  (.D(N_82_i), .CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .EN(N_97_i), .ALn(DB_OUT), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(dly_cnt_Z[0]));
    CFG4 #( .INIT(16'hEEEC) )  \current_state_RNO[12]  (.A(
        current_state_Z[12]), .B(current_state_Z[11]), .C(N_69), .D(
        dly_cnt_Z[4]), .Y(N_284_i));
    CFG2 #( .INIT(4'h8) )  \current_state_RNO[11]  (.A(
        current_state_Z[0]), .B(PLL_LOCK_0), .Y(N_41_i));
    SLE \reset_cycle_count[1]  (.D(N_51_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(reset_cycle_count_Z[1]));
    CFG4 #( .INIT(16'h1000) )  \current_state_ns_a2_1[4]  (.A(
        transition_check_counter_Z[7]), .B(
        transition_check_counter_Z[6]), .C(
        current_state_ns_a2_1_6_Z[4]), .D(current_state_ns_a2_1_5_Z[4])
        , .Y(N_212));
    CFG3 #( .INIT(8'hFB) )  \current_state_ns_0_o2[5]  (.A(
        transition_detected_Z), .B(current_state_Z[5]), .C(
        un1_vcophsel_bclk_1_Z), .Y(N_76));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[0]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[0])
        , .D(GND), .FCI(transition_check_counter_cry_cy), .S(
        transition_check_counter_s[0]), .Y(
        transition_check_counter_cry_Y[0]), .FCO(
        transition_check_counter_cry_Z[0]));
    SLE \bclk_igear_rx_reg[3]  (.D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_374_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        bclk_igear_rx_reg_Z[3]));
    SLE transition_detected (.D(transition_detected_3), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(transition_detected_Z));
    SLE \rotate_count[1]  (.D(N_78_i_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(next_state43_1));
    CFG4 #( .INIT(16'hEEEC) )  \current_state_RNO[10]  (.A(
        current_state_Z[10]), .B(current_state_Z[9]), .C(dly_cnt_Z[4]), 
        .D(N_69), .Y(N_281_i));
    SLE \current_state[8]  (.D(N_38_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[8]));
    CFG3 #( .INIT(8'hFE) )  dly_cnt_n2_i_o2_0 (.A(dly_cnt_Z[2]), .B(
        dly_cnt_Z[1]), .C(dly_cnt_Z[0]), .Y(N_68));
    SLE \current_state[12]  (.D(N_284_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[12]));
    CFG4 #( .INIT(16'h7BDE) )  \register_rx.un4_transition_detected_1  
        (.A(bclk_igear_rx_reg_Z[3]), .B(bclk_igear_rx_reg_Z[2]), .C(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3]), .D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2]), .Y(
        un4_transition_detected_1));
    CFG4 #( .INIT(16'hA9FF) )  dly_cnt_n2_i (.A(dly_cnt_Z[2]), .B(
        dly_cnt_Z[1]), .C(dly_cnt_Z[0]), .D(N_144), .Y(N_23));
    CFG4 #( .INIT(16'hFCEC) )  \current_state_ns_i_a2_i[6]  (.A(
        transition_detected_Z), .B(current_state_Z[8]), .C(
        current_state_Z[5]), .D(un1_vcophsel_bclk_1_Z), .Y(N_64));
    SLE \current_state[1]  (.D(current_state_ns[1]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[1]));
    SLE \current_state[2]  (.D(N_354_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[2]));
    CFG4 #( .INIT(16'hC535) )  \dly_cnt_RNO[4]  (.A(N_62_i), .B(
        dly_cnt_Z[4]), .C(N_144), .D(N_69), .Y(N_91_i));
    SLE \dly_cnt[3]  (.D(N_88_i), .CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .EN(N_97_i), .ALn(DB_OUT), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(dly_cnt_Z[3]));
    CFG4 #( .INIT(16'hEF00) )  \current_state_RNO[8]  (.A(
        next_state43_1), .B(next_state43_0), .C(rotate_count_Z[2]), .D(
        current_state_Z[6]), .Y(N_38_i));
    CFG3 #( .INIT(8'h06) )  \reset_cycle_count_RNO[0]  (.A(
        reset_cycle_count_Z[0]), .B(current_state_Z[4]), .C(
        un1_rst_clk_align_trng_1_0_0_Z), .Y(N_53_i));
    CFG4 #( .INIT(16'h0001) )  \current_state_ns_a2_1_6[4]  (.A(
        transition_check_counter_Z[3]), .B(
        transition_check_counter_Z[2]), .C(
        transition_check_counter_Z[1]), .D(
        transition_check_counter_Z[0]), .Y(
        current_state_ns_a2_1_6_Z[4]));
    CFG4 #( .INIT(16'h0002) )  \current_state_ns_a2_0_a2_0[13]  (.A(
        reset_cycle_count_Z[3]), .B(reset_cycle_count_Z[2]), .C(
        reset_cycle_count_Z[1]), .D(reset_cycle_count_Z[0]), .Y(N_145));
    CFG3 #( .INIT(8'h02) )  \current_state_ns_a2_0_a2[1]  (.A(
        current_state_Z[12]), .B(dly_cnt_Z[4]), .C(N_69), .Y(
        current_state_ns[1]));
    SLE \current_state[4]  (.D(N_59_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[4]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[7]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[7])
        , .D(GND), .FCI(transition_check_counter_cry_Z[6]), .S(
        transition_check_counter_s[7]), .Y(
        transition_check_counter_cry_Y[7]), .FCO(
        transition_check_counter_cry_Z[7]));
    CFG2 #( .INIT(4'hE) )  \current_state_RNIAAGF[8]  (.A(
        current_state_Z[4]), .B(current_state_Z[8]), .Y(N_386_i));
    ARI1 #( .INIT(20'h45500) )  \current_state_RNI00O7[1]  (.A(VCC), 
        .B(current_state_Z[1]), .C(GND), .D(GND), .FCI(VCC), .S(
        current_state_RNI00O7_S[1]), .Y(current_state_RNI00O7_Y_0), 
        .FCO(vcophsel_bclk_cry_cy));
    SLE \current_state[11]  (.D(N_41_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[11]));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNIKA532[2]  (.A(VCC), 
        .B(current_state_Z[1]), .C(vcophsel_bclk_Z[2]), .D(GND), .FCI(
        vcophsel_bclk_cry[1]), .S(vcophsel_bclk_s[2]), .Y(
        vcophsel_bclk_RNIKA532_Y[2]), .FCO(vcophsel_bclk_cry[2]));
    CFG3 #( .INIT(8'h02) )  \current_state_ns_i_0_a2_0[14]  (.A(
        current_state_Z[14]), .B(dly_cnt_Z[4]), .C(N_69), .Y(
        current_state_ns[15]));
    CFG4 #( .INIT(16'hFAF8) )  \current_state_RNO[2]  (.A(
        current_state_Z[2]), .B(dly_cnt_Z[4]), .C(N_126_i), .D(N_69), 
        .Y(N_354_i));
    CFG3 #( .INIT(8'h7F) )  
        \reset_cycle_counter.reset_cycle_count_5_i_o2[2]  (.A(
        reset_cycle_count_Z[1]), .B(reset_cycle_count_Z[0]), .C(
        current_state_Z[4]), .Y(N_72));
    CFG3 #( .INIT(8'hFE) )  \current_state_RNIPT6V[15]  (.A(
        current_state_Z[15]), .B(current_state_Z[1]), .C(
        current_state_Z[5]), .Y(N_374_i));
    SLE \dly_cnt[1]  (.D(N_85_i), .CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .EN(N_97_i), .ALn(DB_OUT), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(dly_cnt_Z[1]));
    CFG2 #( .INIT(4'h1) )  vcophsel_bclk90_sel_0_a2_0_a2 (.A(
        current_state_Z[0]), .B(current_state_0), .Y(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL));
    SLE \current_state[0]  (.D(current_state_ns[0]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[0]));
    SLE \transition_check_counter[3]  (.D(
        transition_check_counter_s[3]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[3]));
    SLE \reset_cycle_count[3]  (.D(N_47_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(reset_cycle_count_Z[3]));
    CFG4 #( .INIT(16'h8880) )  \register_rx.transition_detected_3  (.A(
        un8_transition_detected), .B(un10_transition_detected), .C(
        un4_transition_detected_1), .D(un4_transition_detected_0), .Y(
        transition_detected_3));
    CFG4 #( .INIT(16'hAAAE) )  \current_state_RNO[4]  (.A(
        current_state_Z[15]), .B(N_212), .C(N_145), .D(N_76), .Y(
        N_59_i));
    CFG3 #( .INIT(8'h04) )  \current_state_RNIFOTE1[9]  (.A(
        current_state_Z[4]), .B(N_62_i), .C(current_state_Z[9]), .Y(
        N_144));
    SLE \current_state[14]  (.D(N_287_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[14]));
    ARI1 #( .INIT(20'h42200) )  \transition_check_counter_s[9]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[9])
        , .D(GND), .FCI(transition_check_counter_cry_Z[8]), .S(
        transition_check_counter_s_Z[9]), .Y(
        transition_check_counter_s_Y[9]), .FCO(
        transition_check_counter_s_FCO[9]));
    SLE \vcophsel_bclk[1]  (.D(vcophsel_bclk_s[1]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[1]));
    SLE \transition_check_counter[9]  (.D(
        transition_check_counter_s_Z[9]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[9]));
    SLE \transition_check_counter[5]  (.D(
        transition_check_counter_s[5]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[5]));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNO[6]  (.A(VCC), .B(
        current_state_Z[1]), .C(vcophsel_bclk_Z[6]), .D(GND), .FCI(
        vcophsel_bclk_cry[5]), .S(vcophsel_bclk_s[6]), .Y(
        vcophsel_bclk_RNO_Y[6]), .FCO(vcophsel_bclk_RNO_FCO[6]));
    SLE \transition_check_counter[1]  (.D(
        transition_check_counter_s[1]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[1]));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNIH1PA3[4]  (.A(VCC), 
        .B(current_state_Z[1]), .C(vcophsel_bclk_Z[4]), .D(GND), .FCI(
        vcophsel_bclk_cry[3]), .S(vcophsel_bclk_s[4]), .Y(
        vcophsel_bclk_RNIH1PA3_Y[4]), .FCO(vcophsel_bclk_cry[4]));
    SLE \current_state[15]  (.D(current_state_ns[15]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[15]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[3]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[3])
        , .D(GND), .FCI(transition_check_counter_cry_Z[2]), .S(
        transition_check_counter_s[3]), .Y(
        transition_check_counter_cry_Y[3]), .FCO(
        transition_check_counter_cry_Z[3]));
    SLE \dly_cnt[4]  (.D(N_91_i), .CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .EN(N_97_i), .ALn(DB_OUT), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(dly_cnt_Z[4]));
    CFG3 #( .INIT(8'h6A) )  \rotate_count_RNO[1]  (.A(next_state43_1), 
        .B(next_state43_0), .C(current_state_Z[8]), .Y(N_78_i_i));
    CFG2 #( .INIT(4'h1) )  \dly_cnt_RNINST31[4]  (.A(N_69), .B(
        dly_cnt_Z[4]), .Y(N_315_i_0));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[8]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[8])
        , .D(GND), .FCI(transition_check_counter_cry_Z[7]), .S(
        transition_check_counter_s[8]), .Y(
        transition_check_counter_cry_Y[8]), .FCO(
        transition_check_counter_cry_Z[8]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[1]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[1])
        , .D(GND), .FCI(transition_check_counter_cry_Z[0]), .S(
        transition_check_counter_s[1]), .Y(
        transition_check_counter_cry_Y[1]), .FCO(
        transition_check_counter_cry_Z[1]));
    SLE \transition_check_counter[8]  (.D(
        transition_check_counter_s[8]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[8]));
    SLE \current_state[5]  (.D(current_state_ns[5]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[5]));
    SLE \transition_check_counter[4]  (.D(
        transition_check_counter_s[4]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[4]));
    CFG4 #( .INIT(16'hC535) )  \dly_cnt_RNO[3]  (.A(N_62_i), .B(
        dly_cnt_Z[3]), .C(N_144), .D(N_68), .Y(N_88_i));
    SLE \current_state[6]  (.D(N_64), .CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G)
        , .EN(VCC), .ALn(DB_OUT), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(current_state_Z[6]));
    GND GND_Z (.Y(GND));
    CFG2 #( .INIT(4'hE) )  \current_state_RNI33GF[4]  (.A(
        current_state_Z[1]), .B(current_state_Z[4]), .Y(N_126_i));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'h1000) )  \current_state_ns_a2_0_a2_7[0]  (.A(
        current_state_Z[5]), .B(current_state_Z[8]), .C(
        current_state_ns_a2_0_a2_5_Z[0]), .D(
        current_state_ns_a2_0_a2_3_Z[0]), .Y(
        current_state_ns_a2_0_a2_7_Z[0]));
    SLE \current_state[13]  (.D(current_state_ns[13]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[13]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[2]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[2])
        , .D(GND), .FCI(transition_check_counter_cry_Z[1]), .S(
        transition_check_counter_s[2]), .Y(
        transition_check_counter_cry_Y[2]), .FCO(
        transition_check_counter_cry_Z[2]));
    SLE \transition_check_counter[6]  (.D(
        transition_check_counter_s[6]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(GND)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        transition_check_counter_Z[6]));
    CFG3 #( .INIT(8'h53) )  \dly_cnt_RNO[0]  (.A(dly_cnt_Z[0]), .B(
        N_62_i), .C(N_144), .Y(N_82_i));
    SLE \vcophsel_bclk[4]  (.D(vcophsel_bclk_s[4]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[4]));
    SLE \bclk_igear_rx_reg[2]  (.D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_374_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        bclk_igear_rx_reg_Z[2]));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNINGBF1[1]  (.A(VCC), 
        .B(current_state_Z[1]), .C(vcophsel_bclk_Z[1]), .D(GND), .FCI(
        vcophsel_bclk_cry[0]), .S(vcophsel_bclk_s[1]), .Y(
        vcophsel_bclk_RNINGBF1_Y[1]), .FCO(vcophsel_bclk_cry[1]));
    SLE \current_state[10]  (.D(N_281_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[10]));
    CFG4 #( .INIT(16'h0010) )  un1_vcophsel_bclk_1_4 (.A(
        vcophsel_bclk_Z[5]), .B(vcophsel_bclk_Z[4]), .C(
        vcophsel_bclk_Z[3]), .D(vcophsel_bclk_Z[2]), .Y(
        un1_vcophsel_bclk_1_4_Z));
    CFG4 #( .INIT(16'h0200) )  un1_vcophsel_bclk_1 (.A(
        vcophsel_bclk_Z[6]), .B(vcophsel_bclk_Z[1]), .C(
        vcophsel_bclk_Z[0]), .D(un1_vcophsel_bclk_1_4_Z), .Y(
        un1_vcophsel_bclk_1_Z));
    CFG4 #( .INIT(16'hEEE2) )  \current_state_RNO[14]  (.A(
        current_state_Z[13]), .B(current_state_Z[14]), .C(dly_cnt_Z[4])
        , .D(N_69), .Y(N_287_i));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNIHUIU3[5]  (.A(VCC), 
        .B(current_state_Z[1]), .C(vcophsel_bclk_Z[5]), .D(GND), .FCI(
        vcophsel_bclk_cry[4]), .S(vcophsel_bclk_s[5]), .Y(
        vcophsel_bclk_RNIHUIU3_Y[5]), .FCO(vcophsel_bclk_cry[5]));
    SLE \current_state[7]  (.D(current_state_ns[7]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_0));
    SLE \vcophsel_bclk[5]  (.D(vcophsel_bclk_s[5]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[5]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[6]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[6])
        , .D(GND), .FCI(transition_check_counter_cry_Z[5]), .S(
        transition_check_counter_s[6]), .Y(
        transition_check_counter_cry_Y[6]), .FCO(
        transition_check_counter_cry_Z[6]));
    CFG2 #( .INIT(4'hD) )  reset_lane_i_a3_i_o2 (.A(N_62_i), .B(
        current_state_Z[9]), .Y(N_81));
    SLE \vcophsel_bclk[6]  (.D(vcophsel_bclk_s[6]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[6]));
    CFG3 #( .INIT(8'hEC) )  un1_rst_clk_align_trng_1_0_0 (.A(
        current_state_Z[4]), .B(current_state_Z[1]), .C(N_145), .Y(
        un1_rst_clk_align_trng_1_0_0_Z));
    CFG4 #( .INIT(16'h990F) )  \dly_cnt_RNO[1]  (.A(dly_cnt_Z[1]), .B(
        dly_cnt_Z[0]), .C(N_62_i), .D(N_144), .Y(N_85_i));
    SLE \bclk_igear_rx_reg[1]  (.D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_374_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        bclk_igear_rx_reg_Z[1]));
    CFG4 #( .INIT(16'h6AAA) )  \rotate_count_RNO[2]  (.A(
        rotate_count_Z[2]), .B(next_state43_1), .C(next_state43_0), .D(
        current_state_Z[8]), .Y(rotate_count_4[2]));
    CFG4 #( .INIT(16'h0001) )  \current_state_ns_a2_0_a2_5[0]  (.A(
        current_state_Z[14]), .B(current_state_Z[12]), .C(
        current_state_Z[10]), .D(current_state_Z[6]), .Y(
        current_state_ns_a2_0_a2_5_Z[0]));
    CFG3 #( .INIT(8'h08) )  \current_state_ns_a2_0_a2[13]  (.A(N_212), 
        .B(N_145), .C(N_76), .Y(current_state_ns[13]));
    CFG4 #( .INIT(16'h0002) )  \current_state_ns_a2_0_a2[0]  (.A(
        current_state_ns_a2_0_a2_7_Z[0]), .B(N_81), .C(
        current_state_Z[2]), .D(N_126_i), .Y(current_state_ns[0]));
    CFG2 #( .INIT(4'h1) )  \current_state_RNI4DDV[11]  (.A(
        current_state_Z[11]), .B(current_state_Z[13]), .Y(N_62_i));
    SLE \current_state[9]  (.D(current_state_ns[9]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(current_state_Z[9]));
    ARI1 #( .INIT(20'h44400) )  \vcophsel_bclk_RNII5VM2[3]  (.A(VCC), 
        .B(current_state_Z[1]), .C(vcophsel_bclk_Z[3]), .D(GND), .FCI(
        vcophsel_bclk_cry[2]), .S(vcophsel_bclk_s[3]), .Y(
        vcophsel_bclk_RNII5VM2_Y[3]), .FCO(vcophsel_bclk_cry[3]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[5]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[5])
        , .D(GND), .FCI(transition_check_counter_cry_Z[4]), .S(
        transition_check_counter_s[5]), .Y(
        transition_check_counter_cry_Y[5]), .FCO(
        transition_check_counter_cry_Z[5]));
    ARI1 #( .INIT(20'h62200) )  \transition_check_counter_cry[4]  (.A(
        VCC), .B(current_state_Z[5]), .C(transition_check_counter_Z[4])
        , .D(GND), .FCI(transition_check_counter_cry_Z[3]), .S(
        transition_check_counter_s[4]), .Y(
        transition_check_counter_cry_Y[4]), .FCO(
        transition_check_counter_cry_Z[4]));
    CFG4 #( .INIT(16'h006A) )  \reset_cycle_count_RNO[1]  (.A(
        reset_cycle_count_Z[1]), .B(reset_cycle_count_Z[0]), .C(
        current_state_Z[4]), .D(un1_rst_clk_align_trng_1_0_0_Z), .Y(
        N_51_i));
    SLE \vcophsel_bclk[3]  (.D(vcophsel_bclk_s[3]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_126_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(vcophsel_bclk_Z[3]));
    SLE \reset_cycle_count[0]  (.D(N_53_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(reset_cycle_count_Z[0]));
    CFG4 #( .INIT(16'hEFFF) )  \current_state_RNI6LRI2[9]  (.A(
        current_state_Z[4]), .B(current_state_Z[9]), .C(N_315_i_0), .D(
        N_62_i), .Y(N_97_i));
    CFG4 #( .INIT(16'hECA0) )  \current_state_ns_0[7]  (.A(PLL_LOCK_0), 
        .B(current_state_Z[10]), .C(current_state_0), .D(N_315_i_0), 
        .Y(current_state_ns[7]));
    CFG4 #( .INIT(16'h7BDE) )  \register_rx.un4_transition_detected_0  
        (.A(bclk_igear_rx_reg_Z[1]), .B(bclk_igear_rx_reg_Z[0]), .C(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1]), .D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]), .Y(
        un4_transition_detected_0));
    CFG4 #( .INIT(16'hFFFE) )  \register_rx.un8_transition_detected  (
        .A(PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1]), .B(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]), .C(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3]), .D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2]), .Y(
        un8_transition_detected));
    SLE \bclk_igear_rx_reg[0]  (.D(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(N_374_i), .ALn(DB_OUT), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        bclk_igear_rx_reg_Z[0]));
    SLE \reset_cycle_count[2]  (.D(N_49_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(DB_OUT), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(reset_cycle_count_Z[2]));
    
endmodule


module PF_IOD_TX_CCC_C0_TR_PF_IOD_TX_CCC_C0_TR_0_COREBCLKSCLKALIGN_Z4(
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX,
       current_state_0,
       current_state_RNI00O7_Y_0,
       DB_OUT,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       N_81,
       COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL,
       PLL_LOCK_0,
       N_386_i
    );
input  [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
output current_state_0;
output current_state_RNI00O7_Y_0;
input  DB_OUT;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;
output N_81;
output COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL;
input  PLL_LOCK_0;
output N_386_i;

    wire GND, VCC;
    
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    PLL_BCLKSCLKALIGN_Z5 \genblk1.U_PLL_BCLKSCLKALIGN  (
        .current_state_RNI00O7_Y_0(current_state_RNI00O7_Y_0), 
        .current_state_0(current_state_0), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX({
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]}), .N_386_i(
        N_386_i), .PLL_LOCK_0(PLL_LOCK_0), 
        .COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL), .N_81(N_81), 
        .PF_IOD_TX_CCC_C0_0_TX_CLK_G(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .DB_OUT(DB_OUT));
    
endmodule


module PF_IOD_TX_CCC_C0_TR(
       current_state_RNI00O7_Y_0,
       current_state_0,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX,
       N_386_i,
       PLL_LOCK_0,
       COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL,
       N_81,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       DB_OUT
    );
output current_state_RNI00O7_Y_0;
output current_state_0;
input  [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
output N_386_i;
input  PLL_LOCK_0;
output COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL;
output N_81;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;
input  DB_OUT;

    wire GND, VCC;
    
    PF_IOD_TX_CCC_C0_TR_PF_IOD_TX_CCC_C0_TR_0_COREBCLKSCLKALIGN_Z4 
        PF_IOD_TX_CCC_C0_TR_0 (
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX({
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]}), 
        .current_state_0(current_state_0), .current_state_RNI00O7_Y_0(
        current_state_RNI00O7_Y_0), .DB_OUT(DB_OUT), 
        .PF_IOD_TX_CCC_C0_0_TX_CLK_G(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .N_81(N_81), .COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL), .PLL_LOCK_0(
        PLL_LOCK_0), .N_386_i(N_386_i));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_TX_CCC_C0_PF_CCC_0_PF_CCC(
       current_state_RNI00O7_Y_0,
       PF_CCC_C0_0_OUT0_FABCLK_0,
       COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL,
       N_386_i,
       DB_OUT,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       PLL_LOCK_c_i,
       PLL_LOCK_0,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90
    );
input  current_state_RNI00O7_Y_0;
input  PF_CCC_C0_0_OUT0_FABCLK_0;
input  COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL;
input  N_386_i;
input  DB_OUT;
output PF_IOD_TX_CCC_C0_0_TX_CLK_G;
output PLL_LOCK_c_i;
output PLL_LOCK_0;
output PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0;
output PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90;

    wire [7:0] SSCG_WAVE_TABLE_ADDR;
    wire [32:0] DRI_RDATA;
    wire Y_4, Y_5, pll_inst_0_clkint_8, pll_inst_0_hs_io_clk_3, 
        pll_inst_0_hs_io_clk_7, VCC, GND, DELAY_LINE_OUT_OF_RANGE_1, 
        pll_inst_0_clkint_12, DRI_INTERRUPT;
    
    CLKINT hs_io_clk_7_RNIF7AB (.A(Y_4), .Y(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90));
    CLKINT clkint_8 (.A(pll_inst_0_clkint_8), .Y(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G));
    CFG1 #( .INIT(2'h1) )  pll_inst_0_RNI2EDF (.A(PLL_LOCK_0), .Y(
        PLL_LOCK_c_i));
    PLL #( .VCOFREQUENCY(2000), .DELAY_LINE_SIMULATION_MODE(""), .DATA_RATE(0.000000)
        , .FORMAL_NAME(""), .INTERFACE_NAME(""), .INTERFACE_LEVEL(32'b00000000000000000000000000000000)
        , .SOFTRESET(32'b00000000000000000000000000000000), .SOFT_POWERDOWN_N(32'b00000000000000000000000000000001)
        , .RFDIV_EN(32'b00000000000000000000000000000001), .OUT0_DIV_EN(32'b00000000000000000000000000000001)
        , .OUT1_DIV_EN(32'b00000000000000000000000000000001), .OUT2_DIV_EN(32'b00000000000000000000000000000001)
        , .OUT3_DIV_EN(32'b00000000000000000000000000000001), .SOFT_REF_CLK_SEL(32'b00000000000000000000000000000000)
        , .RESET_ON_LOCK(32'b00000000000000000000000000000001), .BYPASS_CLK_SEL(32'b00000000000000000000000000000000)
        , .BYPASS_GO_EN_N(32'b00000000000000000000000000000001), .BYPASS_PLL(32'b00000000000000000000000000000000)
        , .BYPASS_OUT_DIVIDER(32'b00000000000000000000000000000000), .FF_REQUIRES_LOCK(32'b00000000000000000000000000000000)
        , .FSE_N(32'b00000000000000000000000000000000), .FB_CLK_SEL_0(32'b00000000000000000000000000000000)
        , .FB_CLK_SEL_1(32'b00000000000000000000000000000000), .RFDIV(32'b00000000000000000000000000000001)
        , .FRAC_EN(32'b00000000000000000000000000000000), .FRAC_DAC_EN(32'b00000000000000000000000000000000)
        , .DIV0_RST_DELAY(32'b00000000000000000000000000000000), .DIV0_VAL(32'b00000000000000000000000000000001)
        , .DIV1_RST_DELAY(32'b00000000000000000000000000000000), .DIV1_VAL(32'b00000000000000000000000000000001)
        , .DIV2_RST_DELAY(32'b00000000000000000000000000000000), .DIV2_VAL(32'b00000000000000000000000000000100)
        , .DIV3_RST_DELAY(32'b00000000000000000000000000000000), .DIV3_VAL(32'b00000000000000000000000000000100)
        , .DIV3_CLK_SEL(32'b00000000000000000000000000000000), .BW_INT_CTRL(32'b00000000000000000000000000000000)
        , .BW_PROP_CTRL(32'b00000000000000000000000000000001), .IREF_EN(32'b00000000000000000000000000000001)
        , .IREF_TOGGLE(32'b00000000000000000000000000000000), .LOCK_CNT(32'b00000000000000000000000000001000)
        , .DESKEW_CAL_CNT(32'b00000000000000000000000000000110), .DESKEW_CAL_EN(32'b00000000000000000000000000000001)
        , .DESKEW_CAL_BYPASS(32'b00000000000000000000000000000000), .SYNC_REF_DIV_EN(32'b00000000000000000000000000000000)
        , .SYNC_REF_DIV_EN_2(32'b00000000000000000000000000000000), .OUT0_PHASE_SEL(32'b00000000000000000000000000000000)
        , .OUT1_PHASE_SEL(32'b00000000000000000000000000000010), .OUT2_PHASE_SEL(32'b00000000000000000000000000000000)
        , .OUT3_PHASE_SEL(32'b00000000000000000000000000000000), .SOFT_LOAD_PHASE_N(32'b00000000000000000000000000000001)
        , .SSM_DIV_VAL(32'b00000000000000000000000000000001), .FB_FRAC_VAL(32'b00000000000000000000000000000000)
        , .SSM_SPREAD_MODE(32'b00000000000000000000000000000000), .SSM_MODULATION(32'b00000000000000000000000000000101)
        , .FB_INT_VAL(32'b00000000000000000000000000010000), .SSM_EN_N(32'b00000000000000000000000000000001)
        , .SSM_EXT_WAVE_EN(32'b00000000000000000000000000000000), .SSM_EXT_WAVE_MAX_ADDR(32'b00000000000000000000000000000000)
        , .SSM_RANDOM_EN(32'b00000000000000000000000000000000), .SSM_RANDOM_PATTERN_SEL(32'b00000000000000000000000000000000)
        , .CDMUX0_SEL(32'b00000000000000000000000000000000), .CDMUX1_SEL(32'b00000000000000000000000000000001)
        , .CDMUX2_SEL(32'b00000000000000000000000000000000), .CDELAY0_SEL(32'b00000000000000000000000000000000)
        , .CDELAY0_EN(32'b00000000000000000000000000000000), .DRI_EN(32'b00000000000000000000000000000001)
         )  pll_inst_0 (.LOCK(PLL_LOCK_0), .SSCG_WAVE_TABLE_ADDR({
        SSCG_WAVE_TABLE_ADDR[7], SSCG_WAVE_TABLE_ADDR[6], 
        SSCG_WAVE_TABLE_ADDR[5], SSCG_WAVE_TABLE_ADDR[4], 
        SSCG_WAVE_TABLE_ADDR[3], SSCG_WAVE_TABLE_ADDR[2], 
        SSCG_WAVE_TABLE_ADDR[1], SSCG_WAVE_TABLE_ADDR[0]}), 
        .DELAY_LINE_OUT_OF_RANGE(DELAY_LINE_OUT_OF_RANGE_1), 
        .POWERDOWN_N(DB_OUT), .OUT0_EN(VCC), .OUT1_EN(VCC), .OUT2_EN(
        VCC), .OUT3_EN(VCC), .REF_CLK_SEL(GND), .BYPASS_EN_N(VCC), 
        .LOAD_PHASE_N(current_state_RNI00O7_Y_0), .SSCG_WAVE_TABLE({
        GND, GND, GND, GND, GND, GND, GND, GND}), .PHASE_DIRECTION(VCC)
        , .PHASE_ROTATE(N_386_i), .PHASE_OUT0_SEL(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL), .PHASE_OUT1_SEL(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL), .PHASE_OUT2_SEL(
        GND), .PHASE_OUT3_SEL(GND), .DELAY_LINE_MOVE(GND), 
        .DELAY_LINE_DIRECTION(GND), .DELAY_LINE_WIDE(GND), 
        .DELAY_LINE_LOAD(VCC), .REFCLK_SYNC_EN(GND), .REF_CLK_0(
        PF_CCC_C0_0_OUT0_FABCLK_0), .REF_CLK_1(GND), .FB_CLK(GND), 
        .OUT0(pll_inst_0_hs_io_clk_3), .OUT1(pll_inst_0_hs_io_clk_7), 
        .OUT2(pll_inst_0_clkint_8), .OUT3(pll_inst_0_clkint_12), 
        .DRI_CLK(GND), .DRI_CTRL({GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND}), .DRI_WDATA({GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .DRI_ARST_N(VCC), .DRI_RDATA({DRI_RDATA[32], 
        DRI_RDATA[31], DRI_RDATA[30], DRI_RDATA[29], DRI_RDATA[28], 
        DRI_RDATA[27], DRI_RDATA[26], DRI_RDATA[25], DRI_RDATA[24], 
        DRI_RDATA[23], DRI_RDATA[22], DRI_RDATA[21], DRI_RDATA[20], 
        DRI_RDATA[19], DRI_RDATA[18], DRI_RDATA[17], DRI_RDATA[16], 
        DRI_RDATA[15], DRI_RDATA[14], DRI_RDATA[13], DRI_RDATA[12], 
        DRI_RDATA[11], DRI_RDATA[10], DRI_RDATA[9], DRI_RDATA[8], 
        DRI_RDATA[7], DRI_RDATA[6], DRI_RDATA[5], DRI_RDATA[4], 
        DRI_RDATA[3], DRI_RDATA[2], DRI_RDATA[1], DRI_RDATA[0]}), 
        .DRI_INTERRUPT(DRI_INTERRUPT));
    VCC VCC_Z (.Y(VCC));
    HS_IO_CLK hs_io_clk_7 (.A(pll_inst_0_hs_io_clk_7), .Y(Y_4));
    CLKINT hs_io_clk_3_RNIB7AB (.A(Y_5), .Y(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0));
    HS_IO_CLK hs_io_clk_3 (.A(pll_inst_0_hs_io_clk_3), .Y(Y_5));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_TX_CCC_C0(
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX,
       current_state_0,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0,
       PLL_LOCK_c_i,
       PF_CCC_C0_0_OUT0_FABCLK_0,
       DB_OUT,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       N_81,
       PLL_LOCK_0
    );
input  [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
output current_state_0;
output PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90;
output PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0;
output PLL_LOCK_c_i;
input  PF_CCC_C0_0_OUT0_FABCLK_0;
input  DB_OUT;
output PF_IOD_TX_CCC_C0_0_TX_CLK_G;
output N_81;
output PLL_LOCK_0;

    wire [1:1] current_state_RNI00O7_Y;
    wire N_386_i, COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL, GND, VCC;
    
    PF_IOD_TX_CCC_C0_TR COREBCLKSCLKALIGN_0 (
        .current_state_RNI00O7_Y_0(current_state_RNI00O7_Y[1]), 
        .current_state_0(current_state_0), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX({
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]}), .N_386_i(
        N_386_i), .PLL_LOCK_0(PLL_LOCK_0), 
        .COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL), .N_81(N_81), 
        .PF_IOD_TX_CCC_C0_0_TX_CLK_G(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .DB_OUT(DB_OUT));
    VCC VCC_Z (.Y(VCC));
    PF_IOD_TX_CCC_C0_PF_CCC_0_PF_CCC PF_CCC_0 (
        .current_state_RNI00O7_Y_0(current_state_RNI00O7_Y[1]), 
        .PF_CCC_C0_0_OUT0_FABCLK_0(PF_CCC_C0_0_OUT0_FABCLK_0), 
        .COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL(
        COREBCLKSCLKALIGN_0_PLL_VCOPHSEL_BCLK_SEL), .N_386_i(N_386_i), 
        .DB_OUT(DB_OUT), .PF_IOD_TX_CCC_C0_0_TX_CLK_G(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .PLL_LOCK_c_i(PLL_LOCK_c_i), 
        .PLL_LOCK_0(PLL_LOCK_0), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90));
    GND GND_Z (.Y(GND));
    
endmodule


module ACT_UNIQUE_prbscheck_parallel_fab(
       rev_bits_0_out_data_4,
       PRBS_ERR_0_c,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst
    );
input  [7:0] rev_bits_0_out_data_4;
output PRBS_ERR_0_c;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  RX_CLK_ALIGN_DONE_arst;

    wire [6:0] s_in_old_Z;
    wire [7:0] s_error1_Z;
    wire [0:0] s_error1_2_Z;
    wire [1:1] s_error1_3_Z;
    wire [2:2] s_error1_4_Z;
    wire [3:3] s_error1_5_Z;
    wire [4:4] s_error1_6_Z;
    wire [5:5] s_error1_7_Z;
    wire [6:6] s_error1_8_Z;
    wire [7:7] s_error1_9_Z;
    wire VCC, GND, s_error0_Z, un1_s_error0_i, s_prbs_chk_error_Z, 
        un1_s_error0_4_Z, s_prbs_chk_error_5_Z, s_prbs_chk_error_4_Z;
    
    CFG3 #( .INIT(8'h96) )  \s_error1_8[6]  (.A(s_in_old_Z[4]), .B(
        rev_bits_0_out_data_4[6]), .C(s_in_old_Z[5]), .Y(
        s_error1_8_Z[6]));
    GND GND_Z (.Y(GND));
    SLE \s_in_old[0]  (.D(rev_bits_0_out_data_4[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[0]));
    CFG4 #( .INIT(16'hFFFE) )  un1_s_error0_4 (.A(
        rev_bits_0_out_data_4[3]), .B(rev_bits_0_out_data_4[1]), .C(
        rev_bits_0_out_data_4[2]), .D(rev_bits_0_out_data_4[6]), .Y(
        un1_s_error0_4_Z));
    SLE \s_in_old[6]  (.D(rev_bits_0_out_data_4[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[6]));
    SLE \s_in_old[3]  (.D(rev_bits_0_out_data_4[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[3]));
    SLE \s_error1[7]  (.D(s_error1_9_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[7]));
    VCC VCC_Z (.Y(VCC));
    SLE \s_error1[6]  (.D(s_error1_8_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[6]));
    SLE prbs_chk_error_o (.D(s_prbs_chk_error_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(PRBS_ERR_0_c));
    SLE \s_error1[0]  (.D(s_error1_2_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[0]));
    CFG3 #( .INIT(8'h96) )  \s_error1_6[4]  (.A(s_in_old_Z[2]), .B(
        rev_bits_0_out_data_4[4]), .C(s_in_old_Z[3]), .Y(
        s_error1_6_Z[4]));
    CFG3 #( .INIT(8'h96) )  \s_error1_5[3]  (.A(s_in_old_Z[1]), .B(
        rev_bits_0_out_data_4[3]), .C(s_in_old_Z[2]), .Y(
        s_error1_5_Z[3]));
    SLE \s_error1[1]  (.D(s_error1_3_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[1]));
    CFG4 #( .INIT(16'hFFFE) )  s_prbs_chk_error (.A(s_error1_Z[4]), .B(
        s_error1_Z[5]), .C(s_prbs_chk_error_5_Z), .D(
        s_prbs_chk_error_4_Z), .Y(s_prbs_chk_error_Z));
    SLE \s_in_old[1]  (.D(rev_bits_0_out_data_4[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[1]));
    CFG4 #( .INIT(16'hFFFE) )  s_prbs_chk_error_5 (.A(s_error1_Z[3]), 
        .B(s_error1_Z[2]), .C(s_error1_Z[1]), .D(s_error1_Z[0]), .Y(
        s_prbs_chk_error_5_Z));
    SLE \s_error1[3]  (.D(s_error1_5_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[3]));
    SLE \s_in_old[4]  (.D(rev_bits_0_out_data_4[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[4]));
    CFG3 #( .INIT(8'h96) )  \s_error1_9[7]  (.A(s_in_old_Z[5]), .B(
        rev_bits_0_out_data_4[7]), .C(s_in_old_Z[6]), .Y(
        s_error1_9_Z[7]));
    CFG3 #( .INIT(8'h96) )  \s_error1_2[0]  (.A(
        rev_bits_0_out_data_4[6]), .B(rev_bits_0_out_data_4[7]), .C(
        rev_bits_0_out_data_4[0]), .Y(s_error1_2_Z[0]));
    SLE \s_in_old[5]  (.D(rev_bits_0_out_data_4[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[5]));
    SLE \s_error1[2]  (.D(s_error1_4_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[2]));
    CFG4 #( .INIT(16'h0001) )  s_error0_RNO (.A(
        rev_bits_0_out_data_4[5]), .B(rev_bits_0_out_data_4[0]), .C(
        rev_bits_0_out_data_4[4]), .D(un1_s_error0_4_Z), .Y(
        un1_s_error0_i));
    SLE s_error0 (.D(un1_s_error0_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error0_Z));
    SLE \s_in_old[2]  (.D(rev_bits_0_out_data_4[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[2]));
    CFG3 #( .INIT(8'h96) )  \s_error1_3[1]  (.A(
        rev_bits_0_out_data_4[1]), .B(s_in_old_Z[0]), .C(
        rev_bits_0_out_data_4[7]), .Y(s_error1_3_Z[1]));
    CFG3 #( .INIT(8'h96) )  \s_error1_4[2]  (.A(s_in_old_Z[0]), .B(
        rev_bits_0_out_data_4[2]), .C(s_in_old_Z[1]), .Y(
        s_error1_4_Z[2]));
    CFG3 #( .INIT(8'h96) )  \s_error1_7[5]  (.A(s_in_old_Z[3]), .B(
        rev_bits_0_out_data_4[5]), .C(s_in_old_Z[4]), .Y(
        s_error1_7_Z[5]));
    SLE \s_error1[5]  (.D(s_error1_7_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[5]));
    CFG3 #( .INIT(8'hFE) )  s_prbs_chk_error_4 (.A(s_error1_Z[7]), .B(
        s_error1_Z[6]), .C(s_error0_Z), .Y(s_prbs_chk_error_4_Z));
    SLE \s_error1[4]  (.D(s_error1_6_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[4]));
    
endmodule


module PF_IOD_GENERIC_RX_C1_PF_CLK_DIV_RXCLK_PF_CLK_DIV_DELAY(
       PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK,
       HS_IO_CLK_CASCADED_Y
    );
output PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK;
input  HS_IO_CLK_CASCADED_Y;

    wire GND, VCC, DELAY_LINE_OUT_OF_RANGE, CLK_DIV_OUT, Y_3, Y_ND_0;
    
    ICB_CLKDIVDELAY #( .DELAY_LINE_SIMULATION_MODE("DISABLED"), .DIVIDER(3'b100)
        , .DELAY_LINE_EN(1'b1), .DELAY_LINE_VAL(7'b0000000), .DELAY_VAL_X2(1'b1)
        , .FB_SOURCE_SEL_0(2'b00), .FB_SOURCE_SEL_1(2'b01) )  I_CDD (
        .DELAY_LINE_OUT_OF_RANGE(DELAY_LINE_OUT_OF_RANGE), 
        .DELAY_LINE_DIR(GND), .DELAY_LINE_MOVE(GND), .DELAY_LINE_LOAD(
        GND), .RST_N(VCC), .BIT_SLIP(GND), .A(HS_IO_CLK_CASCADED_Y), 
        .Y_DIV(CLK_DIV_OUT), .Y(Y_3), .Y_FB(
        PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK), .Y_ND(Y_ND_0));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1_PF_CLK_DIV_FIFO_PF_CLK_DIV_DELAY(
       PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK,
       PF_CLK_DIV_FIFO_CLK_DIV_OUT,
       HS_IO_CLK_CASCADED_Y,
       PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV
    );
output PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK;
output PF_CLK_DIV_FIFO_CLK_DIV_OUT;
input  HS_IO_CLK_CASCADED_Y;
output PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE;
input  COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD;
input  COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV;

    wire VCC, GND, Y_2, Y_ND;
    
    ICB_CLKDIVDELAY #( .DELAY_LINE_SIMULATION_MODE("ENABLED"), .DIVIDER(3'b100)
        , .DELAY_LINE_EN(1'b1), .DELAY_LINE_VAL(7'b0000001), .DELAY_VAL_X2(1'b1)
        , .FB_SOURCE_SEL_0(2'b00), .FB_SOURCE_SEL_1(2'b01) )  I_CDD (
        .DELAY_LINE_OUT_OF_RANGE(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), .DELAY_LINE_DIR(VCC), 
        .DELAY_LINE_MOVE(COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV), 
        .DELAY_LINE_LOAD(COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD), 
        .RST_N(VCC), .BIT_SLIP(GND), .A(HS_IO_CLK_CASCADED_Y), .Y_DIV(
        PF_CLK_DIV_FIFO_CLK_DIV_OUT), .Y(Y_2), .Y_FB(
        PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK), .Y_ND(Y_ND));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1_PF_IOD_CLK_TRAINING_PF_IOD(
       PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT,
       HS_IO_CLK_FIFO_Y,
       PF_LANECTRL_0_TX_SYNC_RST,
       PF_LANECTRL_0_RX_SYNC_RST,
       PF_LANECTRL_0_ARST_N,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS
    );
input  [2:0] PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT;
input  HS_IO_CLK_FIFO_Y;
input  PF_LANECTRL_0_TX_SYNC_RST;
input  PF_LANECTRL_0_RX_SYNC_RST;
input  PF_LANECTRL_0_ARST_N;
output PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0;
output PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS;

    wire [1:0] RX_DATA_1;
    wire [9:2] RX_DATA;
    wire [10:0] CDR_CLK_B_SEL_1;
    wire GND, DELAY_LINE_OUT_OF_RANGE_0, TX_1, OE_1, DDR_DO_READ_1, 
        CDR_CLK_A_SEL_8_1, CDR_CLK_A_SEL_9_1, CDR_CLK_A_SEL_10_1, 
        SWITCH_2, CDR_CLR_NEXT_CLK_N_1, TX_DATA_OUT_9_1, 
        TX_DATA_OUT_8_1, AL_N_OUT_1, OUTFF_SL_OUT_1, OUTFF_EN_OUT_1, 
        INFF_SL_OUT_1, INFF_EN_OUT_1, RX_CLK_OUT_1, TX_CLK_OUT_1, VCC;
    
    VCC VCC_Z (.Y(VCC));
    IOD #( .DATA_RATE(500.000000), .FORMAL_NAME("HS_IO_CLK_TRAINING")
        , .INTERFACE_NAME("RX_DDRX_B_G_DYN"), .DELAY_LINE_SIMULATION_MODE("DISABLED")
        , .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000), .RESERVED_0(1'b0)
        , .RX_CLK_EN(1'b1), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b0), .TX_CLK_INV(1'b0)
        , .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b00), .RX_MODE(4'b0100), .EYE_MONITOR_MODE(1'b1)
        , .DYN_DELAY_LINE_EN(1'b0), .FIFO_WR_EN(1'b0), .EYE_MONITOR_EN(1'b1)
        , .TX_MODE(7'b0000000), .TX_CLK_SEL(2'b00), .TX_OE_MODE(3'b111)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b0)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b1)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b11)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_0 (.EYE_MONITOR_EARLY(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), .EYE_MONITOR_LATE(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), .RX_DATA({RX_DATA[9], 
        RX_DATA[8], RX_DATA[7], RX_DATA[6], RX_DATA[5], RX_DATA[4], 
        RX_DATA[3], RX_DATA[2], RX_DATA_1[1], RX_DATA_1[0]}), 
        .DELAY_LINE_OUT_OF_RANGE(DELAY_LINE_OUT_OF_RANGE_0), .TX_DATA({
        GND, GND, GND, GND, GND, GND, GND, GND}), .OE_DATA({GND, GND, 
        GND, GND}), .RX_BIT_SLIP(GND), .EYE_MONITOR_CLEAR_FLAGS(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS), .DELAY_LINE_MOVE(
        GND), .DELAY_LINE_DIRECTION(GND), .DELAY_LINE_LOAD(GND), 
        .RX_CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .TX_CLK(GND), 
        .ODT_EN(GND), .INFF_SL(GND), .INFF_EN(GND), .OUTFF_SL(GND), 
        .OUTFF_EN(GND), .AL_N(GND), .OEFF_LAT_N(GND), .OEFF_SD_N(GND), 
        .OEFF_AD_N(GND), .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(
        GND), .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), 
        .RX_P(GND), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(GND), 
        .ARST_N(PF_LANECTRL_0_ARST_N), .RX_SYNC_RST(
        PF_LANECTRL_0_RX_SYNC_RST), .TX_SYNC_RST(
        PF_LANECTRL_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, GND, 
        GND, HS_IO_CLK_FIFO_Y}), .RX_DQS_90({GND, GND}), .TX_DQS(GND), 
        .TX_DQS_270(GND), .FIFO_WR_PTR({GND, GND, GND}), .FIFO_RD_PTR({
        GND, GND, GND}), .TX(TX_1), .OE(OE_1), .CDR_CLK(GND), 
        .CDR_NEXT_CLK(GND), .EYE_MONITOR_LANE_WIDTH({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), .DDR_DO_READ(
        DDR_DO_READ_1), .CDR_CLK_A_SEL_8(CDR_CLK_A_SEL_8_1), 
        .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9_1), .CDR_CLK_A_SEL_10(
        CDR_CLK_A_SEL_10_1), .CDR_CLK_B_SEL({CDR_CLK_B_SEL_1[10], 
        CDR_CLK_B_SEL_1[9], CDR_CLK_B_SEL_1[8], CDR_CLK_B_SEL_1[7], 
        CDR_CLK_B_SEL_1[6], CDR_CLK_B_SEL_1[5], CDR_CLK_B_SEL_1[4], 
        CDR_CLK_B_SEL_1[3], CDR_CLK_B_SEL_1[2], CDR_CLK_B_SEL_1[1], 
        CDR_CLK_B_SEL_1[0]}), .SWITCH(SWITCH_2), .CDR_CLR_NEXT_CLK_N(
        CDR_CLR_NEXT_CLK_N_1), .TX_DATA_OUT_9(TX_DATA_OUT_9_1), 
        .TX_DATA_OUT_8(TX_DATA_OUT_8_1), .AL_N_OUT(AL_N_OUT_1), 
        .OUTFF_SL_OUT(OUTFF_SL_OUT_1), .OUTFF_EN_OUT(OUTFF_EN_OUT_1), 
        .INFF_SL_OUT(INFF_SL_OUT_1), .INFF_EN_OUT(INFF_EN_OUT_1), 
        .RX_CLK_OUT(RX_CLK_OUT_1), .TX_CLK_OUT(TX_CLK_OUT_1));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1_PF_LANECTRL_0_PF_LANECTRL_PAUSE_SYNC_3(
       current_state_0,
       HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net,
       PAUSE_MX_0_Y,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G
    );
input  current_state_0;
output HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net;
input  PAUSE_MX_0_Y;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;

    wire RX_CLK_G_i, VCC, pause_sync_0_i, GND;
    
    SLE \pipe_fall.pause_sync_0  (.D(PAUSE_MX_0_Y), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(pause_sync_0_i));
    SLE \pipe_fall.pause_sync  (.D(pause_sync_0_i), .CLK(RX_CLK_G_i), 
        .EN(VCC), .ALn(current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND)
        , .LAT(GND), .Q(HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net)
        );
    CFG1 #( .INIT(2'h1) )  \pipe_fall.pause_sync_RNO  (.A(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .Y(RX_CLK_G_i));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1_PF_LANECTRL_0_PF_LANECTRL(
       PF_LANECTRL_0_FIFO_RD_PTR,
       PF_LANECTRL_0_FIFO_WR_PTR,
       PF_LANECTRL_0_RX_DQS_90_0,
       PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT,
       BIT_ALGN_EYE_IN_c,
       current_state_0,
       PAUSE_MX_0_Y,
       PF_LANECTRL_0_TX_SYNC_RST,
       PF_LANECTRL_0_RX_SYNC_RST,
       PF_LANECTRL_0_ARST_N,
       HS_IO_CLK_RX_Y,
       HS_IO_CLK_FIFO_Y,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G
    );
output [2:0] PF_LANECTRL_0_FIFO_RD_PTR;
output [2:0] PF_LANECTRL_0_FIFO_WR_PTR;
output PF_LANECTRL_0_RX_DQS_90_0;
output [2:0] PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT;
input  [2:0] BIT_ALGN_EYE_IN_c;
input  current_state_0;
input  PAUSE_MX_0_Y;
output PF_LANECTRL_0_TX_SYNC_RST;
output PF_LANECTRL_0_RX_SYNC_RST;
output PF_LANECTRL_0_ARST_N;
input  HS_IO_CLK_RX_Y;
input  HS_IO_CLK_FIFO_Y;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;

    wire [1:1] RX_DQS_90;
    wire ARST_N_i, GND, HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net, 
        VCC, RX_DATA_VALID, RX_BURST_DETECT, 
        RX_DELAY_LINE_OUT_OF_RANGE, TX_DELAY_LINE_OUT_OF_RANGE, 
        CLK_OUT_R, A_OUT_RST_N, ODT_EN_SEL, TX_DQS, TX_DQS_270, 
        CDR_CLK, CDR_NEXT_CLK, ODT_EN_OUT;
    
    CFG1 #( .INIT(2'h1) )  I_LANECTRL_RNO (.A(current_state_0), .Y(
        ARST_N_i));
    LANECTRL #( .DATA_RATE(500.000000), .FORMAL_NAME("RX%DUPLICATE"), .INTERFACE_NAME("RX_DDRX_B_G_DYN")
        , .DELAY_LINE_SIMULATION_MODE("DISABLED"), .INTERFACE_LEVEL(3'b000)
        , .RESERVED_0(1'b0), .RESERVED_1(1'b0), .RESERVED_2(1'b0), .SOFTRESET_EN(1'b0)
        , .SOFTRESET(1'b0), .RX_DQS_DELAY_LINE_EN(1'b1), .TX_DQS_DELAY_LINE_EN(1'b0)
        , .RX_DQS_DELAY_LINE_DIRECTION(1'b1), .TX_DQS_DELAY_LINE_DIRECTION(1'b1)
        , .RX_DQS_DELAY_VAL(8'b00000001), .TX_DQS_DELAY_VAL(8'b00000001)
        , .FIFO_EN(1'b1), .FIFO_MODE(1'b0), .FIFO_RD_PTR_MODE(3'b011)
        , .DQS_MODE(3'b011), .CDR_EN(2'b01), .HS_IO_CLK_SEL(9'b111001000)
        , .DLL_CODE_SEL(2'b00), .CDR_CLK_SEL(12'b000000000000), .READ_MARGIN_TEST_EN(1'b1)
        , .WRITE_MARGIN_TEST_EN(1'b0), .CDR_CLK_DIV(3'b100), .DIV_CLK_SEL(2'b00)
        , .HS_IO_CLK_PAUSE_EN(1'b1), .QDR_EN(1'b0), .DYN_ODT_MODE(1'b0)
        , .DIV_CLK_EN_SRC(2'b11), .RANK_2_MODE(1'b0) )  I_LANECTRL (
        .RX_DATA_VALID(RX_DATA_VALID), .RX_BURST_DETECT(
        RX_BURST_DETECT), .RX_DELAY_LINE_OUT_OF_RANGE(
        RX_DELAY_LINE_OUT_OF_RANGE), .TX_DELAY_LINE_OUT_OF_RANGE(
        TX_DELAY_LINE_OUT_OF_RANGE), .CLK_OUT_R(CLK_OUT_R), 
        .A_OUT_RST_N(A_OUT_RST_N), .FAB_CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RESET(ARST_N_i), .DDR_READ(
        GND), .READ_CLK_SEL({GND, GND, GND}), .DELAY_LINE_SEL(GND), 
        .DELAY_LINE_LOAD(GND), .DELAY_LINE_DIRECTION(GND), 
        .DELAY_LINE_MOVE(GND), .HS_IO_CLK_PAUSE(
        HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net), .DIV_CLK_EN_N(
        VCC), .RX_BIT_SLIP(GND), .CDR_CLK_A_SEL({GND, GND, GND, GND, 
        GND, GND, GND, GND}), .EYE_MONITOR_WIDTH_IN({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .ODT_EN(GND), .CODE_UPDATE(GND), .DQS(
        GND), .DQS_N(GND), .HS_IO_CLK({GND, GND, GND, GND, 
        HS_IO_CLK_RX_Y, HS_IO_CLK_FIFO_Y}), .DLL_CODE({GND, GND, GND, 
        GND, GND, GND, GND, GND}), .EYE_MONITOR_WIDTH_OUT({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), .ODT_EN_SEL(
        ODT_EN_SEL), .RX_DQS_90({RX_DQS_90[1], 
        PF_LANECTRL_0_RX_DQS_90_0}), .TX_DQS(TX_DQS), .TX_DQS_270(
        TX_DQS_270), .FIFO_WR_PTR({PF_LANECTRL_0_FIFO_WR_PTR[2], 
        PF_LANECTRL_0_FIFO_WR_PTR[1], PF_LANECTRL_0_FIFO_WR_PTR[0]}), 
        .FIFO_RD_PTR({PF_LANECTRL_0_FIFO_RD_PTR[2], 
        PF_LANECTRL_0_FIFO_RD_PTR[1], PF_LANECTRL_0_FIFO_RD_PTR[0]}), 
        .CDR_CLK(CDR_CLK), .CDR_NEXT_CLK(CDR_NEXT_CLK), .ARST_N(
        PF_LANECTRL_0_ARST_N), .RX_SYNC_RST(PF_LANECTRL_0_RX_SYNC_RST), 
        .TX_SYNC_RST(PF_LANECTRL_0_TX_SYNC_RST), .ODT_EN_OUT(
        ODT_EN_OUT), .DDR_DO_READ(GND), .CDR_CLK_A_SEL_8(GND), 
        .CDR_CLK_A_SEL_9(GND), .CDR_CLK_A_SEL_10(GND), .CDR_CLK_B_SEL({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .SWITCH(GND), .CDR_CLR_NEXT_CLK_N(GND));
    PF_IOD_GENERIC_RX_C1_PF_LANECTRL_0_PF_LANECTRL_PAUSE_SYNC_3 
        I_LANECTRL_PAUSE_SYNC (.current_state_0(current_state_0), 
        .HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net(
        HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net), .PAUSE_MX_0_Y(
        PAUSE_MX_0_Y), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1_PF_IOD_RX_PF_IOD(
       ACT_UNIQUE_rev_bits_0_out_data,
       EYE_MONITOR_LATE_net_0,
       EYE_MONITOR_EARLY_net_0,
       PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT,
       PF_LANECTRL_0_FIFO_RD_PTR,
       PF_LANECTRL_0_FIFO_WR_PTR,
       PF_LANECTRL_0_RX_DQS_90_0,
       rev_bits_0_out_data_4,
       RXD,
       RXD_N,
       BIT_ALGN_OOR_c,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS,
       HS_IO_CLK_FIFO_Y,
       PF_LANECTRL_0_TX_SYNC_RST,
       PF_LANECTRL_0_RX_SYNC_RST,
       PF_LANECTRL_0_ARST_N,
       BIT_ALGN_OOR_0_c,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS
    );
output [7:0] ACT_UNIQUE_rev_bits_0_out_data;
output [1:0] EYE_MONITOR_LATE_net_0;
output [1:0] EYE_MONITOR_EARLY_net_0;
input  [2:0] PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT;
input  [2:0] PF_LANECTRL_0_FIFO_RD_PTR;
input  [2:0] PF_LANECTRL_0_FIFO_WR_PTR;
input  PF_LANECTRL_0_RX_DQS_90_0;
output [7:0] rev_bits_0_out_data_4;
input  [1:0] RXD;
input  [1:0] RXD_N;
output BIT_ALGN_OOR_c;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS;
input  HS_IO_CLK_FIFO_Y;
input  PF_LANECTRL_0_TX_SYNC_RST;
input  PF_LANECTRL_0_RX_SYNC_RST;
input  PF_LANECTRL_0_ARST_N;
output BIT_ALGN_OOR_0_c;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS;

    wire [1:0] RX_DATA;
    wire [10:0] CDR_CLK_B_SEL;
    wire [1:0] RX_DATA_0;
    wire [10:0] CDR_CLK_B_SEL_0;
    wire Y_I_INBUF_DIFF_0_net, Y_I_INBUF_DIFF_1_net, GND, TX, OE, 
        DDR_DO_READ, CDR_CLK_A_SEL_8, CDR_CLK_A_SEL_9, 
        CDR_CLK_A_SEL_10, SWITCH_0, CDR_CLR_NEXT_CLK_N, TX_DATA_OUT_9, 
        TX_DATA_OUT_8, AL_N_OUT, OUTFF_SL_OUT, OUTFF_EN_OUT, 
        INFF_SL_OUT, INFF_EN_OUT, RX_CLK_OUT, TX_CLK_OUT, TX_0, OE_0, 
        DDR_DO_READ_0, CDR_CLK_A_SEL_8_0, CDR_CLK_A_SEL_9_0, 
        CDR_CLK_A_SEL_10_0, SWITCH_1, CDR_CLR_NEXT_CLK_N_0, 
        TX_DATA_OUT_9_0, TX_DATA_OUT_8_0, AL_N_OUT_0, OUTFF_SL_OUT_0, 
        OUTFF_EN_OUT_0, INFF_SL_OUT_0, INFF_EN_OUT_0, RX_CLK_OUT_0, 
        TX_CLK_OUT_0, VCC;
    
    IOD #( .DATA_RATE(500.000000), .FORMAL_NAME("RXD%STATIC_DELAY"), .INTERFACE_NAME("RX_DDRX_B_G_DYN")
        , .DELAY_LINE_SIMULATION_MODE("DISABLED"), .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000)
        , .RESERVED_0(1'b0), .RX_CLK_EN(1'b1), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b0)
        , .TX_CLK_INV(1'b0), .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b01), .RX_MODE(4'b1100), .EYE_MONITOR_MODE(1'b0)
        , .DYN_DELAY_LINE_EN(1'b1), .FIFO_WR_EN(1'b1), .EYE_MONITOR_EN(1'b1)
        , .TX_MODE(7'b0000000), .TX_CLK_SEL(2'b00), .TX_OE_MODE(3'b111)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b1)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b1)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b00)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_1 (.EYE_MONITOR_EARLY(EYE_MONITOR_EARLY_net_0[1]), 
        .EYE_MONITOR_LATE(EYE_MONITOR_LATE_net_0[1]), .RX_DATA({
        ACT_UNIQUE_rev_bits_0_out_data[0], 
        ACT_UNIQUE_rev_bits_0_out_data[1], 
        ACT_UNIQUE_rev_bits_0_out_data[2], 
        ACT_UNIQUE_rev_bits_0_out_data[3], 
        ACT_UNIQUE_rev_bits_0_out_data[4], 
        ACT_UNIQUE_rev_bits_0_out_data[5], 
        ACT_UNIQUE_rev_bits_0_out_data[6], 
        ACT_UNIQUE_rev_bits_0_out_data[7], RX_DATA_0[1], RX_DATA_0[0]})
        , .DELAY_LINE_OUT_OF_RANGE(BIT_ALGN_OOR_c), .TX_DATA({GND, GND, 
        GND, GND, GND, GND, GND, GND}), .OE_DATA({GND, GND, GND, GND}), 
        .RX_BIT_SLIP(GND), .EYE_MONITOR_CLEAR_FLAGS(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS), .DELAY_LINE_MOVE(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE), .DELAY_LINE_DIRECTION(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR), .DELAY_LINE_LOAD(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD), .RX_CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .TX_CLK(GND), .ODT_EN(GND), 
        .INFF_SL(GND), .INFF_EN(GND), .OUTFF_SL(GND), .OUTFF_EN(GND), 
        .AL_N(GND), .OEFF_LAT_N(GND), .OEFF_SD_N(GND), .OEFF_AD_N(GND), 
        .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(GND), 
        .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), .RX_P(
        Y_I_INBUF_DIFF_1_net), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(
        GND), .ARST_N(PF_LANECTRL_0_ARST_N), .RX_SYNC_RST(
        PF_LANECTRL_0_RX_SYNC_RST), .TX_SYNC_RST(
        PF_LANECTRL_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, GND, 
        GND, HS_IO_CLK_FIFO_Y}), .RX_DQS_90({GND, 
        PF_LANECTRL_0_RX_DQS_90_0}), .TX_DQS(GND), .TX_DQS_270(GND), 
        .FIFO_WR_PTR({PF_LANECTRL_0_FIFO_WR_PTR[2], 
        PF_LANECTRL_0_FIFO_WR_PTR[1], PF_LANECTRL_0_FIFO_WR_PTR[0]}), 
        .FIFO_RD_PTR({PF_LANECTRL_0_FIFO_RD_PTR[2], 
        PF_LANECTRL_0_FIFO_RD_PTR[1], PF_LANECTRL_0_FIFO_RD_PTR[0]}), 
        .TX(TX_0), .OE(OE_0), .CDR_CLK(GND), .CDR_NEXT_CLK(GND), 
        .EYE_MONITOR_LANE_WIDTH({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), .DDR_DO_READ(
        DDR_DO_READ_0), .CDR_CLK_A_SEL_8(CDR_CLK_A_SEL_8_0), 
        .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9_0), .CDR_CLK_A_SEL_10(
        CDR_CLK_A_SEL_10_0), .CDR_CLK_B_SEL({CDR_CLK_B_SEL_0[10], 
        CDR_CLK_B_SEL_0[9], CDR_CLK_B_SEL_0[8], CDR_CLK_B_SEL_0[7], 
        CDR_CLK_B_SEL_0[6], CDR_CLK_B_SEL_0[5], CDR_CLK_B_SEL_0[4], 
        CDR_CLK_B_SEL_0[3], CDR_CLK_B_SEL_0[2], CDR_CLK_B_SEL_0[1], 
        CDR_CLK_B_SEL_0[0]}), .SWITCH(SWITCH_1), .CDR_CLR_NEXT_CLK_N(
        CDR_CLR_NEXT_CLK_N_0), .TX_DATA_OUT_9(TX_DATA_OUT_9_0), 
        .TX_DATA_OUT_8(TX_DATA_OUT_8_0), .AL_N_OUT(AL_N_OUT_0), 
        .OUTFF_SL_OUT(OUTFF_SL_OUT_0), .OUTFF_EN_OUT(OUTFF_EN_OUT_0), 
        .INFF_SL_OUT(INFF_SL_OUT_0), .INFF_EN_OUT(INFF_EN_OUT_0), 
        .RX_CLK_OUT(RX_CLK_OUT_0), .TX_CLK_OUT(TX_CLK_OUT_0));
    INBUF_DIFF I_INBUF_DIFF_0 (.PADP(RXD[0]), .PADN(RXD_N[0]), .Y(
        Y_I_INBUF_DIFF_0_net));
    VCC VCC_Z (.Y(VCC));
    IOD #( .DATA_RATE(500.000000), .FORMAL_NAME("RXD:NO_IOD_N_SIDE%STATIC_DELAY")
        , .INTERFACE_NAME("RX_DDRX_B_G_DYN"), .DELAY_LINE_SIMULATION_MODE("DISABLED")
        , .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000), .RESERVED_0(1'b0)
        , .RX_CLK_EN(1'b1), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b0), .TX_CLK_INV(1'b0)
        , .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b01), .RX_MODE(4'b1100), .EYE_MONITOR_MODE(1'b0)
        , .DYN_DELAY_LINE_EN(1'b1), .FIFO_WR_EN(1'b1), .EYE_MONITOR_EN(1'b1)
        , .TX_MODE(7'b0000000), .TX_CLK_SEL(2'b00), .TX_OE_MODE(3'b111)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b1)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b1)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b00)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_0 (.EYE_MONITOR_EARLY(EYE_MONITOR_EARLY_net_0[0]), 
        .EYE_MONITOR_LATE(EYE_MONITOR_LATE_net_0[0]), .RX_DATA({
        rev_bits_0_out_data_4[0], rev_bits_0_out_data_4[1], 
        rev_bits_0_out_data_4[2], rev_bits_0_out_data_4[3], 
        rev_bits_0_out_data_4[4], rev_bits_0_out_data_4[5], 
        rev_bits_0_out_data_4[6], rev_bits_0_out_data_4[7], RX_DATA[1], 
        RX_DATA[0]}), .DELAY_LINE_OUT_OF_RANGE(BIT_ALGN_OOR_0_c), 
        .TX_DATA({GND, GND, GND, GND, GND, GND, GND, GND}), .OE_DATA({
        GND, GND, GND, GND}), .RX_BIT_SLIP(GND), 
        .EYE_MONITOR_CLEAR_FLAGS(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS), .DELAY_LINE_MOVE(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE), .DELAY_LINE_DIRECTION(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR), .DELAY_LINE_LOAD(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD), .RX_CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .TX_CLK(GND), .ODT_EN(GND), 
        .INFF_SL(GND), .INFF_EN(GND), .OUTFF_SL(GND), .OUTFF_EN(GND), 
        .AL_N(GND), .OEFF_LAT_N(GND), .OEFF_SD_N(GND), .OEFF_AD_N(GND), 
        .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(GND), 
        .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), .RX_P(
        Y_I_INBUF_DIFF_0_net), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(
        GND), .ARST_N(PF_LANECTRL_0_ARST_N), .RX_SYNC_RST(
        PF_LANECTRL_0_RX_SYNC_RST), .TX_SYNC_RST(
        PF_LANECTRL_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, GND, 
        GND, HS_IO_CLK_FIFO_Y}), .RX_DQS_90({GND, 
        PF_LANECTRL_0_RX_DQS_90_0}), .TX_DQS(GND), .TX_DQS_270(GND), 
        .FIFO_WR_PTR({PF_LANECTRL_0_FIFO_WR_PTR[2], 
        PF_LANECTRL_0_FIFO_WR_PTR[1], PF_LANECTRL_0_FIFO_WR_PTR[0]}), 
        .FIFO_RD_PTR({PF_LANECTRL_0_FIFO_RD_PTR[2], 
        PF_LANECTRL_0_FIFO_RD_PTR[1], PF_LANECTRL_0_FIFO_RD_PTR[0]}), 
        .TX(TX), .OE(OE), .CDR_CLK(GND), .CDR_NEXT_CLK(GND), 
        .EYE_MONITOR_LANE_WIDTH({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), .DDR_DO_READ(
        DDR_DO_READ), .CDR_CLK_A_SEL_8(CDR_CLK_A_SEL_8), 
        .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9), .CDR_CLK_A_SEL_10(
        CDR_CLK_A_SEL_10), .CDR_CLK_B_SEL({CDR_CLK_B_SEL[10], 
        CDR_CLK_B_SEL[9], CDR_CLK_B_SEL[8], CDR_CLK_B_SEL[7], 
        CDR_CLK_B_SEL[6], CDR_CLK_B_SEL[5], CDR_CLK_B_SEL[4], 
        CDR_CLK_B_SEL[3], CDR_CLK_B_SEL[2], CDR_CLK_B_SEL[1], 
        CDR_CLK_B_SEL[0]}), .SWITCH(SWITCH_0), .CDR_CLR_NEXT_CLK_N(
        CDR_CLR_NEXT_CLK_N), .TX_DATA_OUT_9(TX_DATA_OUT_9), 
        .TX_DATA_OUT_8(TX_DATA_OUT_8), .AL_N_OUT(AL_N_OUT), 
        .OUTFF_SL_OUT(OUTFF_SL_OUT), .OUTFF_EN_OUT(OUTFF_EN_OUT), 
        .INFF_SL_OUT(INFF_SL_OUT), .INFF_EN_OUT(INFF_EN_OUT), 
        .RX_CLK_OUT(RX_CLK_OUT), .TX_CLK_OUT(TX_CLK_OUT));
    INBUF_DIFF I_INBUF_DIFF_1 (.PADP(RXD[1]), .PADN(RXD_N[1]), .Y(
        Y_I_INBUF_DIFF_1_net));
    GND GND_Z (.Y(GND));
    
endmodule


module ICB_BCLKSCLKALIGN_Z3(
       current_state_0,
       PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE,
       PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE,
       CLK_TRAIN_ERROR_c,
       COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0,
       RX_CLK_ALIGN_DONE_arst,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G
    );
input  current_state_0;
input  PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE;
output PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE;
output CLK_TRAIN_ERROR_c;
output COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS;
input  PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0;
input  PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0;
output RX_CLK_ALIGN_DONE_arst;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;

    wire [9:0] rst_cnt_Z;
    wire [8:0] rst_cnt_s;
    wire [7:0] timeout_cnt_Z;
    wire [6:0] timeout_cnt_s;
    wire [7:0] sig_tapcnt_final_1_Z;
    wire [7:0] sig_tapcnt_final_2_Z;
    wire [6:0] sig_tapcnt_final_2_3_Z;
    wire [1:1] cnt_Z;
    wire [127:0] early_flags_msb_Z;
    wire [2:0] wait_cnt_Z;
    wire [2:1] wait_cnt_3;
    wire [6:0] sig_tapcnt_final_1_3_Z;
    wire [127:0] late_flags_lsb_Z;
    wire [127:0] late_flags_msb_Z;
    wire [7:0] early_late_init_val_Z;
    wire [7:0] emflag_cnt_Z;
    wire [7:0] tapcnt_final_Z;
    wire [7:0] tapcnt_final_11;
    wire [7:0] early_late_nxt_val_Z;
    wire [7:0] early_late_start_val_Z;
    wire [127:0] early_flags_lsb_Z;
    wire [7:0] early_late_end_val_Z;
    wire [5:0] clkalign_curr_state_Z;
    wire [5:1] clkalign_curr_state_ns;
    wire [7:0] tapcnt_offset_Z;
    wire [7:0] tapcnt_offset_s;
    wire [7:0] tap_cnt_Z;
    wire [6:0] tap_cnt_s;
    wire [7:7] tap_cnt_s_Z;
    wire [7:7] timeout_cnt_s_Z;
    wire [6:0] emflag_cnt_s;
    wire [7:7] emflag_cnt_s_Z;
    wire [9:9] rst_cnt_s_Z;
    wire [0:0] clkalign_curr_state_RNIJB1J_S;
    wire [0:0] clkalign_curr_state_RNIJB1J_Y;
    wire [6:0] tapcnt_offset_cry;
    wire [0:0] tapcnt_offset_RNIUBO91_Y;
    wire [1:1] tapcnt_offset_RNIADF02_Y;
    wire [2:2] tapcnt_offset_RNINF6N2_Y;
    wire [3:3] tapcnt_offset_RNI5JTD3_Y;
    wire [4:4] tapcnt_offset_RNIKNK44_Y;
    wire [5:5] tapcnt_offset_RNI4TBR4_Y;
    wire [7:7] tapcnt_offset_RNO_FCO;
    wire [7:7] tapcnt_offset_RNO_Y;
    wire [6:6] tapcnt_offset_RNIL33I5_Y;
    wire [0:0] tap_cnt_cry_cy_S;
    wire [0:0] tap_cnt_cry_cy_Y;
    wire [6:0] tap_cnt_cry_Z;
    wire [6:0] tap_cnt_cry_Y;
    wire [7:7] tap_cnt_s_FCO;
    wire [7:7] tap_cnt_s_Y;
    wire [0:0] emflag_cnt_cry_cy_S;
    wire [0:0] emflag_cnt_cry_cy_Y;
    wire [6:0] emflag_cnt_cry_Z;
    wire [6:0] emflag_cnt_cry_Y;
    wire [7:7] emflag_cnt_s_FCO;
    wire [7:7] emflag_cnt_s_Y;
    wire [8:1] rst_cnt_cry_Z;
    wire [8:1] rst_cnt_cry_Y;
    wire [9:9] rst_cnt_s_FCO;
    wire [9:9] rst_cnt_s_Y;
    wire [6:1] timeout_cnt_cry_Z;
    wire [6:1] timeout_cnt_cry_Y;
    wire [7:7] timeout_cnt_s_FCO;
    wire [7:7] timeout_cnt_s_Y;
    wire [0:0] wait_cnt_3_i_0;
    wire [27:27] clkalign_curr_state_d;
    wire [0:0] wait_cnt_3_i_a3_2_0;
    wire [7:0] tapcnt_final_11_iv_0;
    wire [7:0] tapcnt_final_11_iv_1;
    wire RX_CLK_ALIGN_DONE_rep_Z, VCC, RX_CLK_ALIGN_DONE5, GND, CO0_0, 
        CO0_0_i, clkalign_curr_state_s9_0_a3, N_677_i, 
        un3_sig_tapcnt_final_1_cry_7_Z, un2_sig_tapcnt_final_2_cry_7_Z, 
        N_554_i, un1_early_flags_lsb14_i, N_673_i, N_511_i, 
        un1_early_flags_lsb14_1_i, un1_clkalign_curr_state_14_0, 
        un1_clkalign_curr_state_11_0, un1_early_late_nxt_set14_1_0, 
        un1_clkalign_curr_state_15_0, un1_early_late_end_set12_1_0, 
        rx_trng_done_Z, N_2967, un1_clkalign_curr_state_1_0, 
        calc_done_Z, calc_done_0_sqmuxa, un1_clkalign_curr_state_17_0, 
        early_late_end_set_Z, N_515_i, early_late_nxt_set_Z, N_517_i, 
        rx_err_Z, timeout_cnte, N_2939, 
        un1_clkalign_curr_state_0_sqmuxa_8_0, N_2935_i, 
        un1_RX_CLK_ALIGN_LOAD5_0, N_2924_i, 
        un1_clkalign_curr_state_1_sqmuxa_5_0, RX_RESET_LANE5, 
        un1_clkalign_curr_state_0_sqmuxa_3_0, reset_dly_fg_Z, 
        reset_dly_fg4, early_late_start_set_Z, early_late_init_set_Z, 
        clk_align_done_Z, clk_align_start6, un1_internal_rst_en_2_0, 
        N_40_i, early_found_lsb_d_Z, early_found_lsb, 
        late_found_lsb_d_Z, late_found_lsb, early_found_msb_d_Z, 
        early_found_msb, late_found_msb_d_Z, late_found_msb, 
        early_not_found_lsb_d_Z, early_found_lsb_i, 
        late_not_found_lsb_d_Z, late_found_lsb_i, 
        early_not_found_msb_d_Z, early_found_msb_i, 
        late_not_found_msb_d_Z, late_found_msb_i, emflag_cnt_done_d_Z, 
        emflag_cnt_done_Z, tapcnt_final_1_status_Z, 
        sig_tapcnt_final_111_Z, tapcnt_final_2_status_Z, 
        sig_tapcnt_final_210_Z, timeout_fg, 
        early_late_start_end_val_status_Z, 
        early_late_start_end_val_status5, 
        early_late_init_nxt_val_status_Z, 
        early_late_init_nxt_val_status5, start_trng_fg_Z, 
        start_trng_fg6, early_or_late_found_lsb_d_Z, 
        early_or_late_found_lsb_Z, early_or_late_found_msb_d_Z, 
        early_or_late_found_msb_Z, no_early_and_late_found_lsb_d_Z, 
        no_early_and_late_found_lsb_Z, no_early_and_late_found_msb_d_Z, 
        no_early_and_late_found_msb_Z, early_late_start_and_end_set_Z, 
        early_late_start_and_end_set5_Z, early_late_init_and_nxt_set_Z, 
        early_late_init_and_nxt_set5_Z, tapcnt_offsete, tap_cnte, 
        emflag_cnte, tapcnt_offset_cry_cy, tap_cnt_cry_cy, 
        emflag_cnt_cry_cy, N_2979, un2_sig_tapcnt_final_2_cry_0_Z, 
        un2_sig_tapcnt_final_2_cry_0_S, un2_sig_tapcnt_final_2_cry_0_Y, 
        un2_sig_tapcnt_final_2_cry_1_Z, un2_sig_tapcnt_final_2_cry_1_S, 
        un2_sig_tapcnt_final_2_cry_1_Y, un2_sig_tapcnt_final_2_cry_2_Z, 
        un2_sig_tapcnt_final_2_cry_2_S, un2_sig_tapcnt_final_2_cry_2_Y, 
        un2_sig_tapcnt_final_2_cry_3_Z, un2_sig_tapcnt_final_2_cry_3_S, 
        un2_sig_tapcnt_final_2_cry_3_Y, un2_sig_tapcnt_final_2_cry_4_Z, 
        un2_sig_tapcnt_final_2_cry_4_S, un2_sig_tapcnt_final_2_cry_4_Y, 
        un2_sig_tapcnt_final_2_cry_5_Z, un2_sig_tapcnt_final_2_cry_5_S, 
        un2_sig_tapcnt_final_2_cry_5_Y, un2_sig_tapcnt_final_2_cry_6_Z, 
        un2_sig_tapcnt_final_2_cry_6_S, un2_sig_tapcnt_final_2_cry_6_Y, 
        un2_sig_tapcnt_final_2_cry_7_S, un2_sig_tapcnt_final_2_cry_7_Y, 
        un3_sig_tapcnt_final_1_cry_0_Z, un3_sig_tapcnt_final_1_cry_0_S, 
        un3_sig_tapcnt_final_1_cry_0_Y, un3_sig_tapcnt_final_1_cry_1_Z, 
        un3_sig_tapcnt_final_1_cry_1_S, un3_sig_tapcnt_final_1_cry_1_Y, 
        un3_sig_tapcnt_final_1_cry_2_Z, un3_sig_tapcnt_final_1_cry_2_S, 
        un3_sig_tapcnt_final_1_cry_2_Y, un3_sig_tapcnt_final_1_cry_3_Z, 
        un3_sig_tapcnt_final_1_cry_3_S, un3_sig_tapcnt_final_1_cry_3_Y, 
        un3_sig_tapcnt_final_1_cry_4_Z, un3_sig_tapcnt_final_1_cry_4_S, 
        un3_sig_tapcnt_final_1_cry_4_Y, un3_sig_tapcnt_final_1_cry_5_Z, 
        un3_sig_tapcnt_final_1_cry_5_S, un3_sig_tapcnt_final_1_cry_5_Y, 
        un3_sig_tapcnt_final_1_cry_6_Z, un3_sig_tapcnt_final_1_cry_6_S, 
        un3_sig_tapcnt_final_1_cry_6_Y, un3_sig_tapcnt_final_1_cry_7_S, 
        un3_sig_tapcnt_final_1_cry_7_Y, 
        early_late_init_nxt_val_status5_cry_0_Z, 
        early_late_init_nxt_val_status5_cry_0_S, 
        early_late_init_nxt_val_status5_cry_0_Y, 
        early_late_init_nxt_val_status5_cry_1_Z, 
        early_late_init_nxt_val_status5_cry_1_S, 
        early_late_init_nxt_val_status5_cry_1_Y, 
        early_late_init_nxt_val_status5_cry_2_Z, 
        early_late_init_nxt_val_status5_cry_2_S, 
        early_late_init_nxt_val_status5_cry_2_Y, 
        early_late_init_nxt_val_status5_cry_3_Z, 
        early_late_init_nxt_val_status5_cry_3_S, 
        early_late_init_nxt_val_status5_cry_3_Y, 
        early_late_init_nxt_val_status5_cry_4_Z, 
        early_late_init_nxt_val_status5_cry_4_S, 
        early_late_init_nxt_val_status5_cry_4_Y, 
        early_late_init_nxt_val_status5_cry_5_Z, 
        early_late_init_nxt_val_status5_cry_5_S, 
        early_late_init_nxt_val_status5_cry_5_Y, 
        early_late_init_nxt_val_status5_cry_6_Z, 
        early_late_init_nxt_val_status5_cry_6_S, 
        early_late_init_nxt_val_status5_cry_6_Y, 
        early_late_init_nxt_val_status5_cry_7_S, 
        early_late_init_nxt_val_status5_cry_7_Y, 
        early_late_start_end_val_status5_cry_0_Z, 
        early_late_start_end_val_status5_cry_0_S, 
        early_late_start_end_val_status5_cry_0_Y, 
        early_late_start_end_val_status5_cry_1_Z, 
        early_late_start_end_val_status5_cry_1_S, 
        early_late_start_end_val_status5_cry_1_Y, 
        early_late_start_end_val_status5_cry_2_Z, 
        early_late_start_end_val_status5_cry_2_S, 
        early_late_start_end_val_status5_cry_2_Y, 
        early_late_start_end_val_status5_cry_3_Z, 
        early_late_start_end_val_status5_cry_3_S, 
        early_late_start_end_val_status5_cry_3_Y, 
        early_late_start_end_val_status5_cry_4_Z, 
        early_late_start_end_val_status5_cry_4_S, 
        early_late_start_end_val_status5_cry_4_Y, 
        early_late_start_end_val_status5_cry_5_Z, 
        early_late_start_end_val_status5_cry_5_S, 
        early_late_start_end_val_status5_cry_5_Y, 
        early_late_start_end_val_status5_cry_6_Z, 
        early_late_start_end_val_status5_cry_6_S, 
        early_late_start_end_val_status5_cry_6_Y, 
        early_late_start_end_val_status5_cry_7_S, 
        early_late_start_end_val_status5_cry_7_Y, rst_cnt_s_1133_FCO, 
        rst_cnt_s_1133_S, rst_cnt_s_1133_Y, timeout_cnt_s_1134_FCO, 
        timeout_cnt_s_1134_S, timeout_cnt_s_1134_Y, m70_1_0_co1, 
        m70_1_0_wmux_0_S, N_71, N_63, i18_mux, m70_1_0_y0, m70_1_0_co0, 
        m70_1_0_wmux_S, N_46, N_58, early_found_lsb_126_2_1_co1_21, 
        early_found_lsb_126_2_1_wmux_44_S, 
        early_found_lsb_126_2_1_0_y45, early_found_lsb_126_2_1_y3_2, 
        early_found_lsb_126_2_1_y1_2, early_found_lsb_126_2_1_y0_19, 
        early_found_lsb_126_2_1_co0_21, 
        early_found_lsb_126_2_1_wmux_43_S, 
        early_found_lsb_126_2_1_y5_2, early_found_lsb_126_2_1_y7_2, 
        early_found_lsb_126_2_1_co1_20, 
        early_found_lsb_126_2_1_wmux_42_S, 
        early_found_lsb_126_2_1_y0_18, early_found_lsb_126_2_1_co0_20, 
        early_found_lsb_126_2_1_wmux_41_S, 
        early_found_lsb_126_2_1_co1_19, 
        early_found_lsb_126_2_1_wmux_40_S, 
        early_found_lsb_126_2_1_y0_17, early_found_lsb_126_2_1_co0_19, 
        early_found_lsb_126_2_1_wmux_39_S, 
        early_found_lsb_126_2_1_co1_18, 
        early_found_lsb_126_2_1_wmux_38_S, 
        early_found_lsb_126_2_1_y0_16, early_found_lsb_126_2_1_co0_18, 
        early_found_lsb_126_2_1_wmux_37_S, 
        early_found_lsb_126_2_1_co1_17, 
        early_found_lsb_126_2_1_wmux_36_S, 
        early_found_lsb_126_2_1_y0_15, early_found_lsb_126_2_1_co0_17, 
        early_found_lsb_126_2_1_wmux_35_S, 
        early_found_lsb_126_2_1_co1_16, 
        early_found_lsb_126_2_1_wmux_34_S, 
        early_found_lsb_126_2_1_wmux_34_Y, 
        early_found_lsb_126_2_1_co0_16, 
        early_found_lsb_126_2_1_wmux_33_S, 
        early_found_lsb_126_2_1_wmux_33_Y, 
        early_found_lsb_126_2_1_co1_15, 
        early_found_lsb_126_2_1_wmux_32_S, 
        early_found_lsb_126_2_1_0_y33, early_found_lsb_126_2_1_y3_1, 
        early_found_lsb_126_2_1_y1_1, early_found_lsb_126_2_1_y0_14, 
        early_found_lsb_126_2_1_co0_15, 
        early_found_lsb_126_2_1_wmux_31_S, 
        early_found_lsb_126_2_1_y5_1, early_found_lsb_126_2_1_y7_1, 
        early_found_lsb_126_2_1_co1_14, 
        early_found_lsb_126_2_1_wmux_30_S, 
        early_found_lsb_126_2_1_y0_13, early_found_lsb_126_2_1_co0_14, 
        early_found_lsb_126_2_1_wmux_29_S, 
        early_found_lsb_126_2_1_co1_13, 
        early_found_lsb_126_2_1_wmux_28_S, 
        early_found_lsb_126_2_1_y0_12, early_found_lsb_126_2_1_co0_13, 
        early_found_lsb_126_2_1_wmux_27_S, 
        early_found_lsb_126_2_1_co1_12, 
        early_found_lsb_126_2_1_wmux_26_S, 
        early_found_lsb_126_2_1_y0_11, early_found_lsb_126_2_1_co0_12, 
        early_found_lsb_126_2_1_wmux_25_S, 
        early_found_lsb_126_2_1_co1_11, 
        early_found_lsb_126_2_1_wmux_24_S, 
        early_found_lsb_126_2_1_y0_10, early_found_lsb_126_2_1_co0_11, 
        early_found_lsb_126_2_1_wmux_23_S, 
        early_found_lsb_126_2_1_co1_10, 
        early_found_lsb_126_2_1_wmux_22_S, 
        early_found_lsb_126_2_1_wmux_22_Y, 
        early_found_lsb_126_2_1_co0_10, 
        early_found_lsb_126_2_1_wmux_21_S, 
        early_found_lsb_126_2_1_wmux_21_Y, 
        early_found_lsb_126_2_1_co1_9, 
        early_found_lsb_126_2_1_wmux_20_S, 
        early_found_lsb_126_2_1_0_y21, early_found_lsb_126_2_1_y3_0, 
        early_found_lsb_126_2_1_y1_0, early_found_lsb_126_2_1_y0_9, 
        early_found_lsb_126_2_1_co0_9, 
        early_found_lsb_126_2_1_wmux_19_S, 
        early_found_lsb_126_2_1_y5_0, early_found_lsb_126_2_1_y7_0, 
        early_found_lsb_126_2_1_co1_8, 
        early_found_lsb_126_2_1_wmux_18_S, 
        early_found_lsb_126_2_1_y0_8, early_found_lsb_126_2_1_co0_8, 
        early_found_lsb_126_2_1_wmux_17_S, 
        early_found_lsb_126_2_1_co1_7, 
        early_found_lsb_126_2_1_wmux_16_S, 
        early_found_lsb_126_2_1_y0_7, early_found_lsb_126_2_1_co0_7, 
        early_found_lsb_126_2_1_wmux_15_S, 
        early_found_lsb_126_2_1_co1_6, 
        early_found_lsb_126_2_1_wmux_14_S, 
        early_found_lsb_126_2_1_y0_6, early_found_lsb_126_2_1_co0_6, 
        early_found_lsb_126_2_1_wmux_13_S, 
        early_found_lsb_126_2_1_co1_5, 
        early_found_lsb_126_2_1_wmux_12_S, 
        early_found_lsb_126_2_1_y0_5, early_found_lsb_126_2_1_co0_5, 
        early_found_lsb_126_2_1_wmux_11_S, 
        early_found_lsb_126_2_1_co1_4, 
        early_found_lsb_126_2_1_wmux_10_S, 
        early_found_lsb_126_2_1_y0_4, early_found_lsb_126_2_1_0_y9, 
        early_found_lsb_126_2_1_co0_4, 
        early_found_lsb_126_2_1_wmux_9_S, N_1967, 
        early_found_lsb_126_2_1_co1_3, 
        early_found_lsb_126_2_1_wmux_8_S, early_found_lsb_126_2_1_0_y3, 
        early_found_lsb_126_2_1_0_y1, early_found_lsb_126_2_1_y0_3, 
        early_found_lsb_126_2_1_co0_3, 
        early_found_lsb_126_2_1_wmux_7_S, early_found_lsb_126_2_1_0_y5, 
        early_found_lsb_126_2_1_0_y7, early_found_lsb_126_2_1_co1_2, 
        early_found_lsb_126_2_1_wmux_6_S, early_found_lsb_126_2_1_y0_2, 
        early_found_lsb_126_2_1_co0_2, 
        early_found_lsb_126_2_1_wmux_5_S, 
        early_found_lsb_126_2_1_co1_1, 
        early_found_lsb_126_2_1_wmux_4_S, early_found_lsb_126_2_1_y0_1, 
        early_found_lsb_126_2_1_co0_1, 
        early_found_lsb_126_2_1_wmux_3_S, 
        early_found_lsb_126_2_1_co1_0, 
        early_found_lsb_126_2_1_wmux_2_S, early_found_lsb_126_2_1_y0_0, 
        early_found_lsb_126_2_1_co0_0, 
        early_found_lsb_126_2_1_wmux_1_S, 
        early_found_lsb_126_2_1_0_co1, 
        early_found_lsb_126_2_1_wmux_0_S, early_found_lsb_126_2_1_0_y0, 
        early_found_lsb_126_2_1_0_co0, 
        early_found_lsb_126_2_1_0_wmux_S, late_found_lsb_63_2_1_co1_21, 
        late_found_lsb_63_2_1_wmux_44_S, late_found_lsb_63_2_1_0_y45, 
        late_found_lsb_63_2_1_y3_2, late_found_lsb_63_2_1_y1_2, 
        late_found_lsb_63_2_1_y0_19, late_found_lsb_63_2_1_co0_21, 
        late_found_lsb_63_2_1_wmux_43_S, late_found_lsb_63_2_1_y5_2, 
        late_found_lsb_63_2_1_y7_2, late_found_lsb_63_2_1_co1_20, 
        late_found_lsb_63_2_1_wmux_42_S, late_found_lsb_63_2_1_y0_18, 
        late_found_lsb_63_2_1_co0_20, late_found_lsb_63_2_1_wmux_41_S, 
        late_found_lsb_63_2_1_co1_19, late_found_lsb_63_2_1_wmux_40_S, 
        late_found_lsb_63_2_1_y0_17, late_found_lsb_63_2_1_co0_19, 
        late_found_lsb_63_2_1_wmux_39_S, late_found_lsb_63_2_1_co1_18, 
        late_found_lsb_63_2_1_wmux_38_S, late_found_lsb_63_2_1_y0_16, 
        late_found_lsb_63_2_1_co0_18, late_found_lsb_63_2_1_wmux_37_S, 
        late_found_lsb_63_2_1_co1_17, late_found_lsb_63_2_1_wmux_36_S, 
        late_found_lsb_63_2_1_y0_15, late_found_lsb_63_2_1_co0_17, 
        late_found_lsb_63_2_1_wmux_35_S, late_found_lsb_63_2_1_co1_16, 
        late_found_lsb_63_2_1_wmux_34_S, 
        late_found_lsb_63_2_1_wmux_34_Y, late_found_lsb_63_2_1_co0_16, 
        late_found_lsb_63_2_1_wmux_33_S, 
        late_found_lsb_63_2_1_wmux_33_Y, late_found_lsb_63_2_1_co1_15, 
        late_found_lsb_63_2_1_wmux_32_S, late_found_lsb_63_2_1_0_y33, 
        late_found_lsb_63_2_1_y3_1, late_found_lsb_63_2_1_y1_1, 
        late_found_lsb_63_2_1_y0_14, late_found_lsb_63_2_1_co0_15, 
        late_found_lsb_63_2_1_wmux_31_S, late_found_lsb_63_2_1_y5_1, 
        late_found_lsb_63_2_1_y7_1, late_found_lsb_63_2_1_co1_14, 
        late_found_lsb_63_2_1_wmux_30_S, late_found_lsb_63_2_1_y0_13, 
        late_found_lsb_63_2_1_co0_14, late_found_lsb_63_2_1_wmux_29_S, 
        late_found_lsb_63_2_1_co1_13, late_found_lsb_63_2_1_wmux_28_S, 
        late_found_lsb_63_2_1_y0_12, late_found_lsb_63_2_1_co0_13, 
        late_found_lsb_63_2_1_wmux_27_S, late_found_lsb_63_2_1_co1_12, 
        late_found_lsb_63_2_1_wmux_26_S, late_found_lsb_63_2_1_y0_11, 
        late_found_lsb_63_2_1_co0_12, late_found_lsb_63_2_1_wmux_25_S, 
        late_found_lsb_63_2_1_co1_11, late_found_lsb_63_2_1_wmux_24_S, 
        late_found_lsb_63_2_1_y0_10, late_found_lsb_63_2_1_co0_11, 
        late_found_lsb_63_2_1_wmux_23_S, late_found_lsb_63_2_1_co1_10, 
        late_found_lsb_63_2_1_wmux_22_S, 
        late_found_lsb_63_2_1_wmux_22_Y, late_found_lsb_63_2_1_co0_10, 
        late_found_lsb_63_2_1_wmux_21_S, 
        late_found_lsb_63_2_1_wmux_21_Y, late_found_lsb_63_2_1_co1_9, 
        late_found_lsb_63_2_1_wmux_20_S, late_found_lsb_63_2_1_0_y21, 
        late_found_lsb_63_2_1_y3_0, late_found_lsb_63_2_1_y1_0, 
        late_found_lsb_63_2_1_y0_9, late_found_lsb_63_2_1_co0_9, 
        late_found_lsb_63_2_1_wmux_19_S, late_found_lsb_63_2_1_y5_0, 
        late_found_lsb_63_2_1_y7_0, late_found_lsb_63_2_1_co1_8, 
        late_found_lsb_63_2_1_wmux_18_S, late_found_lsb_63_2_1_y0_8, 
        late_found_lsb_63_2_1_co0_8, late_found_lsb_63_2_1_wmux_17_S, 
        late_found_lsb_63_2_1_co1_7, late_found_lsb_63_2_1_wmux_16_S, 
        late_found_lsb_63_2_1_y0_7, late_found_lsb_63_2_1_co0_7, 
        late_found_lsb_63_2_1_wmux_15_S, late_found_lsb_63_2_1_co1_6, 
        late_found_lsb_63_2_1_wmux_14_S, late_found_lsb_63_2_1_y0_6, 
        late_found_lsb_63_2_1_co0_6, late_found_lsb_63_2_1_wmux_13_S, 
        late_found_lsb_63_2_1_co1_5, late_found_lsb_63_2_1_wmux_12_S, 
        late_found_lsb_63_2_1_y0_5, late_found_lsb_63_2_1_co0_5, 
        late_found_lsb_63_2_1_wmux_11_S, late_found_lsb_63_2_1_co1_4, 
        late_found_lsb_63_2_1_wmux_10_S, late_found_lsb_63_2_1_y0_4, 
        late_found_lsb_63_2_1_0_y9, late_found_lsb_63_2_1_co0_4, 
        late_found_lsb_63_2_1_wmux_9_S, N_2031, 
        late_found_lsb_63_2_1_co1_3, late_found_lsb_63_2_1_wmux_8_S, 
        late_found_lsb_63_2_1_0_y3, late_found_lsb_63_2_1_0_y1, 
        late_found_lsb_63_2_1_y0_3, late_found_lsb_63_2_1_co0_3, 
        late_found_lsb_63_2_1_wmux_7_S, late_found_lsb_63_2_1_0_y5, 
        late_found_lsb_63_2_1_0_y7, late_found_lsb_63_2_1_co1_2, 
        late_found_lsb_63_2_1_wmux_6_S, late_found_lsb_63_2_1_y0_2, 
        late_found_lsb_63_2_1_co0_2, late_found_lsb_63_2_1_wmux_5_S, 
        late_found_lsb_63_2_1_co1_1, late_found_lsb_63_2_1_wmux_4_S, 
        late_found_lsb_63_2_1_y0_1, late_found_lsb_63_2_1_co0_1, 
        late_found_lsb_63_2_1_wmux_3_S, late_found_lsb_63_2_1_co1_0, 
        late_found_lsb_63_2_1_wmux_2_S, late_found_lsb_63_2_1_y0_0, 
        late_found_lsb_63_2_1_co0_0, late_found_lsb_63_2_1_wmux_1_S, 
        late_found_lsb_63_2_1_0_co1, late_found_lsb_63_2_1_wmux_0_S, 
        late_found_lsb_63_2_1_0_y0, late_found_lsb_63_2_1_0_co0, 
        late_found_lsb_63_2_1_0_wmux_S, early_found_msb_63_2_1_co1_21, 
        early_found_msb_63_2_1_wmux_44_S, early_found_msb_63_2_1_0_y45, 
        early_found_msb_63_2_1_y3_2, early_found_msb_63_2_1_y1_2, 
        early_found_msb_63_2_1_y0_19, early_found_msb_63_2_1_co0_21, 
        early_found_msb_63_2_1_wmux_43_S, early_found_msb_63_2_1_y5_2, 
        early_found_msb_63_2_1_y7_2, early_found_msb_63_2_1_co1_20, 
        early_found_msb_63_2_1_wmux_42_S, early_found_msb_63_2_1_y0_18, 
        early_found_msb_63_2_1_co0_20, 
        early_found_msb_63_2_1_wmux_41_S, 
        early_found_msb_63_2_1_co1_19, 
        early_found_msb_63_2_1_wmux_40_S, early_found_msb_63_2_1_y0_17, 
        early_found_msb_63_2_1_co0_19, 
        early_found_msb_63_2_1_wmux_39_S, 
        early_found_msb_63_2_1_co1_18, 
        early_found_msb_63_2_1_wmux_38_S, early_found_msb_63_2_1_y0_16, 
        early_found_msb_63_2_1_co0_18, 
        early_found_msb_63_2_1_wmux_37_S, 
        early_found_msb_63_2_1_co1_17, 
        early_found_msb_63_2_1_wmux_36_S, early_found_msb_63_2_1_y0_15, 
        early_found_msb_63_2_1_co0_17, 
        early_found_msb_63_2_1_wmux_35_S, 
        early_found_msb_63_2_1_co1_16, 
        early_found_msb_63_2_1_wmux_34_S, 
        early_found_msb_63_2_1_wmux_34_Y, 
        early_found_msb_63_2_1_co0_16, 
        early_found_msb_63_2_1_wmux_33_S, 
        early_found_msb_63_2_1_wmux_33_Y, 
        early_found_msb_63_2_1_co1_15, 
        early_found_msb_63_2_1_wmux_32_S, early_found_msb_63_2_1_0_y33, 
        early_found_msb_63_2_1_y3_1, early_found_msb_63_2_1_y1_1, 
        early_found_msb_63_2_1_y0_14, early_found_msb_63_2_1_co0_15, 
        early_found_msb_63_2_1_wmux_31_S, early_found_msb_63_2_1_y5_1, 
        early_found_msb_63_2_1_y7_1, early_found_msb_63_2_1_co1_14, 
        early_found_msb_63_2_1_wmux_30_S, early_found_msb_63_2_1_y0_13, 
        early_found_msb_63_2_1_co0_14, 
        early_found_msb_63_2_1_wmux_29_S, 
        early_found_msb_63_2_1_co1_13, 
        early_found_msb_63_2_1_wmux_28_S, early_found_msb_63_2_1_y0_12, 
        early_found_msb_63_2_1_co0_13, 
        early_found_msb_63_2_1_wmux_27_S, 
        early_found_msb_63_2_1_co1_12, 
        early_found_msb_63_2_1_wmux_26_S, early_found_msb_63_2_1_y0_11, 
        early_found_msb_63_2_1_co0_12, 
        early_found_msb_63_2_1_wmux_25_S, 
        early_found_msb_63_2_1_co1_11, 
        early_found_msb_63_2_1_wmux_24_S, early_found_msb_63_2_1_y0_10, 
        early_found_msb_63_2_1_co0_11, 
        early_found_msb_63_2_1_wmux_23_S, 
        early_found_msb_63_2_1_co1_10, 
        early_found_msb_63_2_1_wmux_22_S, 
        early_found_msb_63_2_1_wmux_22_Y, 
        early_found_msb_63_2_1_co0_10, 
        early_found_msb_63_2_1_wmux_21_S, 
        early_found_msb_63_2_1_wmux_21_Y, early_found_msb_63_2_1_co1_9, 
        early_found_msb_63_2_1_wmux_20_S, early_found_msb_63_2_1_0_y21, 
        early_found_msb_63_2_1_y3_0, early_found_msb_63_2_1_y1_0, 
        early_found_msb_63_2_1_y0_9, early_found_msb_63_2_1_co0_9, 
        early_found_msb_63_2_1_wmux_19_S, early_found_msb_63_2_1_y5_0, 
        early_found_msb_63_2_1_y7_0, early_found_msb_63_2_1_co1_8, 
        early_found_msb_63_2_1_wmux_18_S, early_found_msb_63_2_1_y0_8, 
        early_found_msb_63_2_1_co0_8, early_found_msb_63_2_1_wmux_17_S, 
        early_found_msb_63_2_1_co1_7, early_found_msb_63_2_1_wmux_16_S, 
        early_found_msb_63_2_1_y0_7, early_found_msb_63_2_1_co0_7, 
        early_found_msb_63_2_1_wmux_15_S, early_found_msb_63_2_1_co1_6, 
        early_found_msb_63_2_1_wmux_14_S, early_found_msb_63_2_1_y0_6, 
        early_found_msb_63_2_1_co0_6, early_found_msb_63_2_1_wmux_13_S, 
        early_found_msb_63_2_1_co1_5, early_found_msb_63_2_1_wmux_12_S, 
        early_found_msb_63_2_1_y0_5, early_found_msb_63_2_1_co0_5, 
        early_found_msb_63_2_1_wmux_11_S, early_found_msb_63_2_1_co1_4, 
        early_found_msb_63_2_1_wmux_10_S, early_found_msb_63_2_1_y0_4, 
        early_found_msb_63_2_1_0_y9, early_found_msb_63_2_1_co0_4, 
        early_found_msb_63_2_1_wmux_9_S, N_2158, 
        early_found_msb_63_2_1_co1_3, early_found_msb_63_2_1_wmux_8_S, 
        early_found_msb_63_2_1_0_y3, early_found_msb_63_2_1_0_y1, 
        early_found_msb_63_2_1_y0_3, early_found_msb_63_2_1_co0_3, 
        early_found_msb_63_2_1_wmux_7_S, early_found_msb_63_2_1_0_y5, 
        early_found_msb_63_2_1_0_y7, early_found_msb_63_2_1_co1_2, 
        early_found_msb_63_2_1_wmux_6_S, early_found_msb_63_2_1_y0_2, 
        early_found_msb_63_2_1_co0_2, early_found_msb_63_2_1_wmux_5_S, 
        early_found_msb_63_2_1_co1_1, early_found_msb_63_2_1_wmux_4_S, 
        early_found_msb_63_2_1_y0_1, early_found_msb_63_2_1_co0_1, 
        early_found_msb_63_2_1_wmux_3_S, early_found_msb_63_2_1_co1_0, 
        early_found_msb_63_2_1_wmux_2_S, early_found_msb_63_2_1_y0_0, 
        early_found_msb_63_2_1_co0_0, early_found_msb_63_2_1_wmux_1_S, 
        early_found_msb_63_2_1_0_co1, early_found_msb_63_2_1_wmux_0_S, 
        early_found_msb_63_2_1_0_y0, early_found_msb_63_2_1_0_co0, 
        early_found_msb_63_2_1_0_wmux_S, 
        early_found_msb_126_2_1_co1_21, 
        early_found_msb_126_2_1_wmux_44_S, 
        early_found_msb_126_2_1_0_y45, early_found_msb_126_2_1_y3_2, 
        early_found_msb_126_2_1_y1_2, early_found_msb_126_2_1_y0_19, 
        early_found_msb_126_2_1_co0_21, 
        early_found_msb_126_2_1_wmux_43_S, 
        early_found_msb_126_2_1_y5_2, early_found_msb_126_2_1_y7_2, 
        early_found_msb_126_2_1_co1_20, 
        early_found_msb_126_2_1_wmux_42_S, 
        early_found_msb_126_2_1_y0_18, early_found_msb_126_2_1_co0_20, 
        early_found_msb_126_2_1_wmux_41_S, 
        early_found_msb_126_2_1_co1_19, 
        early_found_msb_126_2_1_wmux_40_S, 
        early_found_msb_126_2_1_y0_17, early_found_msb_126_2_1_co0_19, 
        early_found_msb_126_2_1_wmux_39_S, 
        early_found_msb_126_2_1_co1_18, 
        early_found_msb_126_2_1_wmux_38_S, 
        early_found_msb_126_2_1_y0_16, early_found_msb_126_2_1_co0_18, 
        early_found_msb_126_2_1_wmux_37_S, 
        early_found_msb_126_2_1_co1_17, 
        early_found_msb_126_2_1_wmux_36_S, 
        early_found_msb_126_2_1_y0_15, early_found_msb_126_2_1_co0_17, 
        early_found_msb_126_2_1_wmux_35_S, 
        early_found_msb_126_2_1_co1_16, 
        early_found_msb_126_2_1_wmux_34_S, 
        early_found_msb_126_2_1_wmux_34_Y, 
        early_found_msb_126_2_1_co0_16, 
        early_found_msb_126_2_1_wmux_33_S, 
        early_found_msb_126_2_1_wmux_33_Y, 
        early_found_msb_126_2_1_co1_15, 
        early_found_msb_126_2_1_wmux_32_S, 
        early_found_msb_126_2_1_0_y33, early_found_msb_126_2_1_y3_1, 
        early_found_msb_126_2_1_y1_1, early_found_msb_126_2_1_y0_14, 
        early_found_msb_126_2_1_co0_15, 
        early_found_msb_126_2_1_wmux_31_S, 
        early_found_msb_126_2_1_y5_1, early_found_msb_126_2_1_y7_1, 
        early_found_msb_126_2_1_co1_14, 
        early_found_msb_126_2_1_wmux_30_S, 
        early_found_msb_126_2_1_y0_13, early_found_msb_126_2_1_co0_14, 
        early_found_msb_126_2_1_wmux_29_S, 
        early_found_msb_126_2_1_co1_13, 
        early_found_msb_126_2_1_wmux_28_S, 
        early_found_msb_126_2_1_y0_12, early_found_msb_126_2_1_co0_13, 
        early_found_msb_126_2_1_wmux_27_S, 
        early_found_msb_126_2_1_co1_12, 
        early_found_msb_126_2_1_wmux_26_S, 
        early_found_msb_126_2_1_y0_11, early_found_msb_126_2_1_co0_12, 
        early_found_msb_126_2_1_wmux_25_S, 
        early_found_msb_126_2_1_co1_11, 
        early_found_msb_126_2_1_wmux_24_S, 
        early_found_msb_126_2_1_y0_10, early_found_msb_126_2_1_co0_11, 
        early_found_msb_126_2_1_wmux_23_S, 
        early_found_msb_126_2_1_co1_10, 
        early_found_msb_126_2_1_wmux_22_S, 
        early_found_msb_126_2_1_wmux_22_Y, 
        early_found_msb_126_2_1_co0_10, 
        early_found_msb_126_2_1_wmux_21_S, 
        early_found_msb_126_2_1_wmux_21_Y, 
        early_found_msb_126_2_1_co1_9, 
        early_found_msb_126_2_1_wmux_20_S, 
        early_found_msb_126_2_1_0_y21, early_found_msb_126_2_1_y3_0, 
        early_found_msb_126_2_1_y1_0, early_found_msb_126_2_1_y0_9, 
        early_found_msb_126_2_1_co0_9, 
        early_found_msb_126_2_1_wmux_19_S, 
        early_found_msb_126_2_1_y5_0, early_found_msb_126_2_1_y7_0, 
        early_found_msb_126_2_1_co1_8, 
        early_found_msb_126_2_1_wmux_18_S, 
        early_found_msb_126_2_1_y0_8, early_found_msb_126_2_1_co0_8, 
        early_found_msb_126_2_1_wmux_17_S, 
        early_found_msb_126_2_1_co1_7, 
        early_found_msb_126_2_1_wmux_16_S, 
        early_found_msb_126_2_1_y0_7, early_found_msb_126_2_1_co0_7, 
        early_found_msb_126_2_1_wmux_15_S, 
        early_found_msb_126_2_1_co1_6, 
        early_found_msb_126_2_1_wmux_14_S, 
        early_found_msb_126_2_1_y0_6, early_found_msb_126_2_1_co0_6, 
        early_found_msb_126_2_1_wmux_13_S, 
        early_found_msb_126_2_1_co1_5, 
        early_found_msb_126_2_1_wmux_12_S, 
        early_found_msb_126_2_1_y0_5, early_found_msb_126_2_1_co0_5, 
        early_found_msb_126_2_1_wmux_11_S, 
        early_found_msb_126_2_1_co1_4, 
        early_found_msb_126_2_1_wmux_10_S, 
        early_found_msb_126_2_1_y0_4, early_found_msb_126_2_1_0_y9, 
        early_found_msb_126_2_1_co0_4, 
        early_found_msb_126_2_1_wmux_9_S, N_2221, 
        early_found_msb_126_2_1_co1_3, 
        early_found_msb_126_2_1_wmux_8_S, early_found_msb_126_2_1_0_y3, 
        early_found_msb_126_2_1_0_y1, early_found_msb_126_2_1_y0_3, 
        early_found_msb_126_2_1_co0_3, 
        early_found_msb_126_2_1_wmux_7_S, early_found_msb_126_2_1_0_y5, 
        early_found_msb_126_2_1_0_y7, early_found_msb_126_2_1_co1_2, 
        early_found_msb_126_2_1_wmux_6_S, early_found_msb_126_2_1_y0_2, 
        early_found_msb_126_2_1_co0_2, 
        early_found_msb_126_2_1_wmux_5_S, 
        early_found_msb_126_2_1_co1_1, 
        early_found_msb_126_2_1_wmux_4_S, early_found_msb_126_2_1_y0_1, 
        early_found_msb_126_2_1_co0_1, 
        early_found_msb_126_2_1_wmux_3_S, 
        early_found_msb_126_2_1_co1_0, 
        early_found_msb_126_2_1_wmux_2_S, early_found_msb_126_2_1_y0_0, 
        early_found_msb_126_2_1_co0_0, 
        early_found_msb_126_2_1_wmux_1_S, 
        early_found_msb_126_2_1_0_co1, 
        early_found_msb_126_2_1_wmux_0_S, early_found_msb_126_2_1_0_y0, 
        early_found_msb_126_2_1_0_co0, 
        early_found_msb_126_2_1_0_wmux_S, late_found_msb_63_2_1_co1_21, 
        late_found_msb_63_2_1_wmux_44_S, late_found_msb_63_2_1_0_y45, 
        late_found_msb_63_2_1_y3_2, late_found_msb_63_2_1_y1_2, 
        late_found_msb_63_2_1_y0_19, late_found_msb_63_2_1_co0_21, 
        late_found_msb_63_2_1_wmux_43_S, late_found_msb_63_2_1_y5_2, 
        late_found_msb_63_2_1_y7_2, late_found_msb_63_2_1_co1_20, 
        late_found_msb_63_2_1_wmux_42_S, late_found_msb_63_2_1_y0_18, 
        late_found_msb_63_2_1_co0_20, late_found_msb_63_2_1_wmux_41_S, 
        late_found_msb_63_2_1_co1_19, late_found_msb_63_2_1_wmux_40_S, 
        late_found_msb_63_2_1_y0_17, late_found_msb_63_2_1_co0_19, 
        late_found_msb_63_2_1_wmux_39_S, late_found_msb_63_2_1_co1_18, 
        late_found_msb_63_2_1_wmux_38_S, late_found_msb_63_2_1_y0_16, 
        late_found_msb_63_2_1_co0_18, late_found_msb_63_2_1_wmux_37_S, 
        late_found_msb_63_2_1_co1_17, late_found_msb_63_2_1_wmux_36_S, 
        late_found_msb_63_2_1_y0_15, late_found_msb_63_2_1_co0_17, 
        late_found_msb_63_2_1_wmux_35_S, late_found_msb_63_2_1_co1_16, 
        late_found_msb_63_2_1_wmux_34_S, 
        late_found_msb_63_2_1_wmux_34_Y, late_found_msb_63_2_1_co0_16, 
        late_found_msb_63_2_1_wmux_33_S, 
        late_found_msb_63_2_1_wmux_33_Y, late_found_msb_63_2_1_co1_15, 
        late_found_msb_63_2_1_wmux_32_S, late_found_msb_63_2_1_0_y33, 
        late_found_msb_63_2_1_y3_1, late_found_msb_63_2_1_y1_1, 
        late_found_msb_63_2_1_y0_14, late_found_msb_63_2_1_co0_15, 
        late_found_msb_63_2_1_wmux_31_S, late_found_msb_63_2_1_y5_1, 
        late_found_msb_63_2_1_y7_1, late_found_msb_63_2_1_co1_14, 
        late_found_msb_63_2_1_wmux_30_S, late_found_msb_63_2_1_y0_13, 
        late_found_msb_63_2_1_co0_14, late_found_msb_63_2_1_wmux_29_S, 
        late_found_msb_63_2_1_co1_13, late_found_msb_63_2_1_wmux_28_S, 
        late_found_msb_63_2_1_y0_12, late_found_msb_63_2_1_co0_13, 
        late_found_msb_63_2_1_wmux_27_S, late_found_msb_63_2_1_co1_12, 
        late_found_msb_63_2_1_wmux_26_S, late_found_msb_63_2_1_y0_11, 
        late_found_msb_63_2_1_co0_12, late_found_msb_63_2_1_wmux_25_S, 
        late_found_msb_63_2_1_co1_11, late_found_msb_63_2_1_wmux_24_S, 
        late_found_msb_63_2_1_y0_10, late_found_msb_63_2_1_co0_11, 
        late_found_msb_63_2_1_wmux_23_S, late_found_msb_63_2_1_co1_10, 
        late_found_msb_63_2_1_wmux_22_S, 
        late_found_msb_63_2_1_wmux_22_Y, late_found_msb_63_2_1_co0_10, 
        late_found_msb_63_2_1_wmux_21_S, 
        late_found_msb_63_2_1_wmux_21_Y, late_found_msb_63_2_1_co1_9, 
        late_found_msb_63_2_1_wmux_20_S, late_found_msb_63_2_1_0_y21, 
        late_found_msb_63_2_1_y3_0, late_found_msb_63_2_1_y1_0, 
        late_found_msb_63_2_1_y0_9, late_found_msb_63_2_1_co0_9, 
        late_found_msb_63_2_1_wmux_19_S, late_found_msb_63_2_1_y5_0, 
        late_found_msb_63_2_1_y7_0, late_found_msb_63_2_1_co1_8, 
        late_found_msb_63_2_1_wmux_18_S, late_found_msb_63_2_1_y0_8, 
        late_found_msb_63_2_1_co0_8, late_found_msb_63_2_1_wmux_17_S, 
        late_found_msb_63_2_1_co1_7, late_found_msb_63_2_1_wmux_16_S, 
        late_found_msb_63_2_1_y0_7, late_found_msb_63_2_1_co0_7, 
        late_found_msb_63_2_1_wmux_15_S, late_found_msb_63_2_1_co1_6, 
        late_found_msb_63_2_1_wmux_14_S, late_found_msb_63_2_1_y0_6, 
        late_found_msb_63_2_1_co0_6, late_found_msb_63_2_1_wmux_13_S, 
        late_found_msb_63_2_1_co1_5, late_found_msb_63_2_1_wmux_12_S, 
        late_found_msb_63_2_1_y0_5, late_found_msb_63_2_1_co0_5, 
        late_found_msb_63_2_1_wmux_11_S, late_found_msb_63_2_1_co1_4, 
        late_found_msb_63_2_1_wmux_10_S, late_found_msb_63_2_1_y0_4, 
        late_found_msb_63_2_1_0_y9, late_found_msb_63_2_1_co0_4, 
        late_found_msb_63_2_1_wmux_9_S, N_2285, 
        late_found_msb_63_2_1_co1_3, late_found_msb_63_2_1_wmux_8_S, 
        late_found_msb_63_2_1_0_y3, late_found_msb_63_2_1_0_y1, 
        late_found_msb_63_2_1_y0_3, late_found_msb_63_2_1_co0_3, 
        late_found_msb_63_2_1_wmux_7_S, late_found_msb_63_2_1_0_y5, 
        late_found_msb_63_2_1_0_y7, late_found_msb_63_2_1_co1_2, 
        late_found_msb_63_2_1_wmux_6_S, late_found_msb_63_2_1_y0_2, 
        late_found_msb_63_2_1_co0_2, late_found_msb_63_2_1_wmux_5_S, 
        late_found_msb_63_2_1_co1_1, late_found_msb_63_2_1_wmux_4_S, 
        late_found_msb_63_2_1_y0_1, late_found_msb_63_2_1_co0_1, 
        late_found_msb_63_2_1_wmux_3_S, late_found_msb_63_2_1_co1_0, 
        late_found_msb_63_2_1_wmux_2_S, late_found_msb_63_2_1_y0_0, 
        late_found_msb_63_2_1_co0_0, late_found_msb_63_2_1_wmux_1_S, 
        late_found_msb_63_2_1_0_co1, late_found_msb_63_2_1_wmux_0_S, 
        late_found_msb_63_2_1_0_y0, late_found_msb_63_2_1_0_co0, 
        late_found_msb_63_2_1_0_wmux_S, late_found_msb_126_2_1_co1_21, 
        late_found_msb_126_2_1_wmux_44_S, late_found_msb_126_2_1_0_y45, 
        late_found_msb_126_2_1_y3_2, late_found_msb_126_2_1_y1_2, 
        late_found_msb_126_2_1_y0_19, late_found_msb_126_2_1_co0_21, 
        late_found_msb_126_2_1_wmux_43_S, late_found_msb_126_2_1_y5_2, 
        late_found_msb_126_2_1_y7_2, late_found_msb_126_2_1_co1_20, 
        late_found_msb_126_2_1_wmux_42_S, late_found_msb_126_2_1_y0_18, 
        late_found_msb_126_2_1_co0_20, 
        late_found_msb_126_2_1_wmux_41_S, 
        late_found_msb_126_2_1_co1_19, 
        late_found_msb_126_2_1_wmux_40_S, late_found_msb_126_2_1_y0_17, 
        late_found_msb_126_2_1_co0_19, 
        late_found_msb_126_2_1_wmux_39_S, 
        late_found_msb_126_2_1_co1_18, 
        late_found_msb_126_2_1_wmux_38_S, late_found_msb_126_2_1_y0_16, 
        late_found_msb_126_2_1_co0_18, 
        late_found_msb_126_2_1_wmux_37_S, 
        late_found_msb_126_2_1_co1_17, 
        late_found_msb_126_2_1_wmux_36_S, late_found_msb_126_2_1_y0_15, 
        late_found_msb_126_2_1_co0_17, 
        late_found_msb_126_2_1_wmux_35_S, 
        late_found_msb_126_2_1_co1_16, 
        late_found_msb_126_2_1_wmux_34_S, 
        late_found_msb_126_2_1_wmux_34_Y, 
        late_found_msb_126_2_1_co0_16, 
        late_found_msb_126_2_1_wmux_33_S, 
        late_found_msb_126_2_1_wmux_33_Y, 
        late_found_msb_126_2_1_co1_15, 
        late_found_msb_126_2_1_wmux_32_S, late_found_msb_126_2_1_0_y33, 
        late_found_msb_126_2_1_y3_1, late_found_msb_126_2_1_y1_1, 
        late_found_msb_126_2_1_y0_14, late_found_msb_126_2_1_co0_15, 
        late_found_msb_126_2_1_wmux_31_S, late_found_msb_126_2_1_y5_1, 
        late_found_msb_126_2_1_y7_1, late_found_msb_126_2_1_co1_14, 
        late_found_msb_126_2_1_wmux_30_S, late_found_msb_126_2_1_y0_13, 
        late_found_msb_126_2_1_co0_14, 
        late_found_msb_126_2_1_wmux_29_S, 
        late_found_msb_126_2_1_co1_13, 
        late_found_msb_126_2_1_wmux_28_S, late_found_msb_126_2_1_y0_12, 
        late_found_msb_126_2_1_co0_13, 
        late_found_msb_126_2_1_wmux_27_S, 
        late_found_msb_126_2_1_co1_12, 
        late_found_msb_126_2_1_wmux_26_S, late_found_msb_126_2_1_y0_11, 
        late_found_msb_126_2_1_co0_12, 
        late_found_msb_126_2_1_wmux_25_S, 
        late_found_msb_126_2_1_co1_11, 
        late_found_msb_126_2_1_wmux_24_S, late_found_msb_126_2_1_y0_10, 
        late_found_msb_126_2_1_co0_11, 
        late_found_msb_126_2_1_wmux_23_S, 
        late_found_msb_126_2_1_co1_10, 
        late_found_msb_126_2_1_wmux_22_S, 
        late_found_msb_126_2_1_wmux_22_Y, 
        late_found_msb_126_2_1_co0_10, 
        late_found_msb_126_2_1_wmux_21_S, 
        late_found_msb_126_2_1_wmux_21_Y, late_found_msb_126_2_1_co1_9, 
        late_found_msb_126_2_1_wmux_20_S, late_found_msb_126_2_1_0_y21, 
        late_found_msb_126_2_1_y3_0, late_found_msb_126_2_1_y1_0, 
        late_found_msb_126_2_1_y0_9, late_found_msb_126_2_1_co0_9, 
        late_found_msb_126_2_1_wmux_19_S, late_found_msb_126_2_1_y5_0, 
        late_found_msb_126_2_1_y7_0, late_found_msb_126_2_1_co1_8, 
        late_found_msb_126_2_1_wmux_18_S, late_found_msb_126_2_1_y0_8, 
        late_found_msb_126_2_1_co0_8, late_found_msb_126_2_1_wmux_17_S, 
        late_found_msb_126_2_1_co1_7, late_found_msb_126_2_1_wmux_16_S, 
        late_found_msb_126_2_1_y0_7, late_found_msb_126_2_1_co0_7, 
        late_found_msb_126_2_1_wmux_15_S, late_found_msb_126_2_1_co1_6, 
        late_found_msb_126_2_1_wmux_14_S, late_found_msb_126_2_1_y0_6, 
        late_found_msb_126_2_1_co0_6, late_found_msb_126_2_1_wmux_13_S, 
        late_found_msb_126_2_1_co1_5, late_found_msb_126_2_1_wmux_12_S, 
        late_found_msb_126_2_1_y0_5, late_found_msb_126_2_1_co0_5, 
        late_found_msb_126_2_1_wmux_11_S, late_found_msb_126_2_1_co1_4, 
        late_found_msb_126_2_1_wmux_10_S, late_found_msb_126_2_1_y0_4, 
        late_found_msb_126_2_1_0_y9, late_found_msb_126_2_1_co0_4, 
        late_found_msb_126_2_1_wmux_9_S, N_2348, 
        late_found_msb_126_2_1_co1_3, late_found_msb_126_2_1_wmux_8_S, 
        late_found_msb_126_2_1_0_y3, late_found_msb_126_2_1_0_y1, 
        late_found_msb_126_2_1_y0_3, late_found_msb_126_2_1_co0_3, 
        late_found_msb_126_2_1_wmux_7_S, late_found_msb_126_2_1_0_y5, 
        late_found_msb_126_2_1_0_y7, late_found_msb_126_2_1_co1_2, 
        late_found_msb_126_2_1_wmux_6_S, late_found_msb_126_2_1_y0_2, 
        late_found_msb_126_2_1_co0_2, late_found_msb_126_2_1_wmux_5_S, 
        late_found_msb_126_2_1_co1_1, late_found_msb_126_2_1_wmux_4_S, 
        late_found_msb_126_2_1_y0_1, late_found_msb_126_2_1_co0_1, 
        late_found_msb_126_2_1_wmux_3_S, late_found_msb_126_2_1_co1_0, 
        late_found_msb_126_2_1_wmux_2_S, late_found_msb_126_2_1_y0_0, 
        late_found_msb_126_2_1_co0_0, late_found_msb_126_2_1_wmux_1_S, 
        late_found_msb_126_2_1_0_co1, late_found_msb_126_2_1_wmux_0_S, 
        late_found_msb_126_2_1_0_y0, late_found_msb_126_2_1_0_co0, 
        late_found_msb_126_2_1_0_wmux_S, late_found_lsb_126_2_1_co1_21, 
        late_found_lsb_126_2_1_wmux_44_S, late_found_lsb_126_2_1_0_y45, 
        late_found_lsb_126_2_1_y3_2, late_found_lsb_126_2_1_y1_2, 
        late_found_lsb_126_2_1_y0_19, late_found_lsb_126_2_1_co0_21, 
        late_found_lsb_126_2_1_wmux_43_S, late_found_lsb_126_2_1_y5_2, 
        late_found_lsb_126_2_1_y7_2, late_found_lsb_126_2_1_co1_20, 
        late_found_lsb_126_2_1_wmux_42_S, late_found_lsb_126_2_1_y0_18, 
        late_found_lsb_126_2_1_co0_20, 
        late_found_lsb_126_2_1_wmux_41_S, 
        late_found_lsb_126_2_1_co1_19, 
        late_found_lsb_126_2_1_wmux_40_S, late_found_lsb_126_2_1_y0_17, 
        late_found_lsb_126_2_1_co0_19, 
        late_found_lsb_126_2_1_wmux_39_S, 
        late_found_lsb_126_2_1_co1_18, 
        late_found_lsb_126_2_1_wmux_38_S, late_found_lsb_126_2_1_y0_16, 
        late_found_lsb_126_2_1_co0_18, 
        late_found_lsb_126_2_1_wmux_37_S, 
        late_found_lsb_126_2_1_co1_17, 
        late_found_lsb_126_2_1_wmux_36_S, late_found_lsb_126_2_1_y0_15, 
        late_found_lsb_126_2_1_co0_17, 
        late_found_lsb_126_2_1_wmux_35_S, 
        late_found_lsb_126_2_1_co1_16, 
        late_found_lsb_126_2_1_wmux_34_S, 
        late_found_lsb_126_2_1_wmux_34_Y, 
        late_found_lsb_126_2_1_co0_16, 
        late_found_lsb_126_2_1_wmux_33_S, 
        late_found_lsb_126_2_1_wmux_33_Y, 
        late_found_lsb_126_2_1_co1_15, 
        late_found_lsb_126_2_1_wmux_32_S, late_found_lsb_126_2_1_0_y33, 
        late_found_lsb_126_2_1_y3_1, late_found_lsb_126_2_1_y1_1, 
        late_found_lsb_126_2_1_y0_14, late_found_lsb_126_2_1_co0_15, 
        late_found_lsb_126_2_1_wmux_31_S, late_found_lsb_126_2_1_y5_1, 
        late_found_lsb_126_2_1_y7_1, late_found_lsb_126_2_1_co1_14, 
        late_found_lsb_126_2_1_wmux_30_S, late_found_lsb_126_2_1_y0_13, 
        late_found_lsb_126_2_1_co0_14, 
        late_found_lsb_126_2_1_wmux_29_S, 
        late_found_lsb_126_2_1_co1_13, 
        late_found_lsb_126_2_1_wmux_28_S, late_found_lsb_126_2_1_y0_12, 
        late_found_lsb_126_2_1_co0_13, 
        late_found_lsb_126_2_1_wmux_27_S, 
        late_found_lsb_126_2_1_co1_12, 
        late_found_lsb_126_2_1_wmux_26_S, late_found_lsb_126_2_1_y0_11, 
        late_found_lsb_126_2_1_co0_12, 
        late_found_lsb_126_2_1_wmux_25_S, 
        late_found_lsb_126_2_1_co1_11, 
        late_found_lsb_126_2_1_wmux_24_S, late_found_lsb_126_2_1_y0_10, 
        late_found_lsb_126_2_1_co0_11, 
        late_found_lsb_126_2_1_wmux_23_S, 
        late_found_lsb_126_2_1_co1_10, 
        late_found_lsb_126_2_1_wmux_22_S, 
        late_found_lsb_126_2_1_wmux_22_Y, 
        late_found_lsb_126_2_1_co0_10, 
        late_found_lsb_126_2_1_wmux_21_S, 
        late_found_lsb_126_2_1_wmux_21_Y, late_found_lsb_126_2_1_co1_9, 
        late_found_lsb_126_2_1_wmux_20_S, late_found_lsb_126_2_1_0_y21, 
        late_found_lsb_126_2_1_y3_0, late_found_lsb_126_2_1_y1_0, 
        late_found_lsb_126_2_1_y0_9, late_found_lsb_126_2_1_co0_9, 
        late_found_lsb_126_2_1_wmux_19_S, late_found_lsb_126_2_1_y5_0, 
        late_found_lsb_126_2_1_y7_0, late_found_lsb_126_2_1_co1_8, 
        late_found_lsb_126_2_1_wmux_18_S, late_found_lsb_126_2_1_y0_8, 
        late_found_lsb_126_2_1_co0_8, late_found_lsb_126_2_1_wmux_17_S, 
        late_found_lsb_126_2_1_co1_7, late_found_lsb_126_2_1_wmux_16_S, 
        late_found_lsb_126_2_1_y0_7, late_found_lsb_126_2_1_co0_7, 
        late_found_lsb_126_2_1_wmux_15_S, late_found_lsb_126_2_1_co1_6, 
        late_found_lsb_126_2_1_wmux_14_S, late_found_lsb_126_2_1_y0_6, 
        late_found_lsb_126_2_1_co0_6, late_found_lsb_126_2_1_wmux_13_S, 
        late_found_lsb_126_2_1_co1_5, late_found_lsb_126_2_1_wmux_12_S, 
        late_found_lsb_126_2_1_y0_5, late_found_lsb_126_2_1_co0_5, 
        late_found_lsb_126_2_1_wmux_11_S, late_found_lsb_126_2_1_co1_4, 
        late_found_lsb_126_2_1_wmux_10_S, late_found_lsb_126_2_1_y0_4, 
        late_found_lsb_126_2_1_0_y9, late_found_lsb_126_2_1_co0_4, 
        late_found_lsb_126_2_1_wmux_9_S, N_2094, 
        late_found_lsb_126_2_1_co1_3, late_found_lsb_126_2_1_wmux_8_S, 
        late_found_lsb_126_2_1_0_y3, late_found_lsb_126_2_1_0_y1, 
        late_found_lsb_126_2_1_y0_3, late_found_lsb_126_2_1_co0_3, 
        late_found_lsb_126_2_1_wmux_7_S, late_found_lsb_126_2_1_0_y5, 
        late_found_lsb_126_2_1_0_y7, late_found_lsb_126_2_1_co1_2, 
        late_found_lsb_126_2_1_wmux_6_S, late_found_lsb_126_2_1_y0_2, 
        late_found_lsb_126_2_1_co0_2, late_found_lsb_126_2_1_wmux_5_S, 
        late_found_lsb_126_2_1_co1_1, late_found_lsb_126_2_1_wmux_4_S, 
        late_found_lsb_126_2_1_y0_1, late_found_lsb_126_2_1_co0_1, 
        late_found_lsb_126_2_1_wmux_3_S, late_found_lsb_126_2_1_co1_0, 
        late_found_lsb_126_2_1_wmux_2_S, late_found_lsb_126_2_1_y0_0, 
        late_found_lsb_126_2_1_co0_0, late_found_lsb_126_2_1_wmux_1_S, 
        late_found_lsb_126_2_1_0_co1, late_found_lsb_126_2_1_wmux_0_S, 
        late_found_lsb_126_2_1_0_y0, late_found_lsb_126_2_1_0_co0, 
        late_found_lsb_126_2_1_0_wmux_S, early_found_lsb_63_2_1_co1_21, 
        early_found_lsb_63_2_1_wmux_44_S, early_found_lsb_63_2_1_0_y45, 
        early_found_lsb_63_2_1_y3_2, early_found_lsb_63_2_1_y1_2, 
        early_found_lsb_63_2_1_y0_19, early_found_lsb_63_2_1_co0_21, 
        early_found_lsb_63_2_1_wmux_43_S, early_found_lsb_63_2_1_y5_2, 
        early_found_lsb_63_2_1_y7_2, early_found_lsb_63_2_1_co1_20, 
        early_found_lsb_63_2_1_wmux_42_S, early_found_lsb_63_2_1_y0_18, 
        early_found_lsb_63_2_1_co0_20, 
        early_found_lsb_63_2_1_wmux_41_S, 
        early_found_lsb_63_2_1_co1_19, 
        early_found_lsb_63_2_1_wmux_40_S, early_found_lsb_63_2_1_y0_17, 
        early_found_lsb_63_2_1_co0_19, 
        early_found_lsb_63_2_1_wmux_39_S, 
        early_found_lsb_63_2_1_co1_18, 
        early_found_lsb_63_2_1_wmux_38_S, early_found_lsb_63_2_1_y0_16, 
        early_found_lsb_63_2_1_co0_18, 
        early_found_lsb_63_2_1_wmux_37_S, 
        early_found_lsb_63_2_1_co1_17, 
        early_found_lsb_63_2_1_wmux_36_S, early_found_lsb_63_2_1_y0_15, 
        early_found_lsb_63_2_1_co0_17, 
        early_found_lsb_63_2_1_wmux_35_S, 
        early_found_lsb_63_2_1_co1_16, 
        early_found_lsb_63_2_1_wmux_34_S, 
        early_found_lsb_63_2_1_wmux_34_Y, 
        early_found_lsb_63_2_1_co0_16, 
        early_found_lsb_63_2_1_wmux_33_S, 
        early_found_lsb_63_2_1_wmux_33_Y, 
        early_found_lsb_63_2_1_co1_15, 
        early_found_lsb_63_2_1_wmux_32_S, early_found_lsb_63_2_1_0_y33, 
        early_found_lsb_63_2_1_y3_1, early_found_lsb_63_2_1_y1_1, 
        early_found_lsb_63_2_1_y0_14, early_found_lsb_63_2_1_co0_15, 
        early_found_lsb_63_2_1_wmux_31_S, early_found_lsb_63_2_1_y5_1, 
        early_found_lsb_63_2_1_y7_1, early_found_lsb_63_2_1_co1_14, 
        early_found_lsb_63_2_1_wmux_30_S, early_found_lsb_63_2_1_y0_13, 
        early_found_lsb_63_2_1_co0_14, 
        early_found_lsb_63_2_1_wmux_29_S, 
        early_found_lsb_63_2_1_co1_13, 
        early_found_lsb_63_2_1_wmux_28_S, early_found_lsb_63_2_1_y0_12, 
        early_found_lsb_63_2_1_co0_13, 
        early_found_lsb_63_2_1_wmux_27_S, 
        early_found_lsb_63_2_1_co1_12, 
        early_found_lsb_63_2_1_wmux_26_S, early_found_lsb_63_2_1_y0_11, 
        early_found_lsb_63_2_1_co0_12, 
        early_found_lsb_63_2_1_wmux_25_S, 
        early_found_lsb_63_2_1_co1_11, 
        early_found_lsb_63_2_1_wmux_24_S, early_found_lsb_63_2_1_y0_10, 
        early_found_lsb_63_2_1_co0_11, 
        early_found_lsb_63_2_1_wmux_23_S, 
        early_found_lsb_63_2_1_co1_10, 
        early_found_lsb_63_2_1_wmux_22_S, 
        early_found_lsb_63_2_1_wmux_22_Y, 
        early_found_lsb_63_2_1_co0_10, 
        early_found_lsb_63_2_1_wmux_21_S, 
        early_found_lsb_63_2_1_wmux_21_Y, early_found_lsb_63_2_1_co1_9, 
        early_found_lsb_63_2_1_wmux_20_S, early_found_lsb_63_2_1_0_y21, 
        early_found_lsb_63_2_1_y3_0, early_found_lsb_63_2_1_y1_0, 
        early_found_lsb_63_2_1_y0_9, early_found_lsb_63_2_1_co0_9, 
        early_found_lsb_63_2_1_wmux_19_S, early_found_lsb_63_2_1_y5_0, 
        early_found_lsb_63_2_1_y7_0, early_found_lsb_63_2_1_co1_8, 
        early_found_lsb_63_2_1_wmux_18_S, early_found_lsb_63_2_1_y0_8, 
        early_found_lsb_63_2_1_co0_8, early_found_lsb_63_2_1_wmux_17_S, 
        early_found_lsb_63_2_1_co1_7, early_found_lsb_63_2_1_wmux_16_S, 
        early_found_lsb_63_2_1_y0_7, early_found_lsb_63_2_1_co0_7, 
        early_found_lsb_63_2_1_wmux_15_S, early_found_lsb_63_2_1_co1_6, 
        early_found_lsb_63_2_1_wmux_14_S, early_found_lsb_63_2_1_y0_6, 
        early_found_lsb_63_2_1_co0_6, early_found_lsb_63_2_1_wmux_13_S, 
        early_found_lsb_63_2_1_co1_5, early_found_lsb_63_2_1_wmux_12_S, 
        early_found_lsb_63_2_1_y0_5, early_found_lsb_63_2_1_co0_5, 
        early_found_lsb_63_2_1_wmux_11_S, early_found_lsb_63_2_1_co1_4, 
        early_found_lsb_63_2_1_wmux_10_S, early_found_lsb_63_2_1_y0_4, 
        early_found_lsb_63_2_1_0_y9, early_found_lsb_63_2_1_co0_4, 
        early_found_lsb_63_2_1_wmux_9_S, N_1904, 
        early_found_lsb_63_2_1_co1_3, early_found_lsb_63_2_1_wmux_8_S, 
        early_found_lsb_63_2_1_0_y3, early_found_lsb_63_2_1_0_y1, 
        early_found_lsb_63_2_1_y0_3, early_found_lsb_63_2_1_co0_3, 
        early_found_lsb_63_2_1_wmux_7_S, early_found_lsb_63_2_1_0_y5, 
        early_found_lsb_63_2_1_0_y7, early_found_lsb_63_2_1_co1_2, 
        early_found_lsb_63_2_1_wmux_6_S, early_found_lsb_63_2_1_y0_2, 
        early_found_lsb_63_2_1_co0_2, early_found_lsb_63_2_1_wmux_5_S, 
        early_found_lsb_63_2_1_co1_1, early_found_lsb_63_2_1_wmux_4_S, 
        early_found_lsb_63_2_1_y0_1, early_found_lsb_63_2_1_co0_1, 
        early_found_lsb_63_2_1_wmux_3_S, early_found_lsb_63_2_1_co1_0, 
        early_found_lsb_63_2_1_wmux_2_S, early_found_lsb_63_2_1_y0_0, 
        early_found_lsb_63_2_1_co0_0, early_found_lsb_63_2_1_wmux_1_S, 
        early_found_lsb_63_2_1_0_co1, early_found_lsb_63_2_1_wmux_0_S, 
        early_found_lsb_63_2_1_0_y0, early_found_lsb_63_2_1_0_co0, 
        early_found_lsb_63_2_1_0_wmux_S, N_643, N_526, N_642, 
        un1_clkalign_curr_state_0_sqmuxa_8_0_0, N_525, N_533, 
        early_or_late_found_Z, N_109, N_61, N_627, N_78, N_546, N_540, 
        N_32_i, N_4, m37_2_1_1_0, N_511_i_1, N_537, m104_1_2, N_97, 
        N_105, N_102, N_82_i, m86_1_0, m86_2, N_87, N_19_i, m57_1_2, 
        N_55, N_130_mux, m74_1_0, N_75, N_30, m54_1_2, m96_1_0, 
        N_139_mux, m114_2_1, N_115, N_137_mux, N_12, m16_2_0_1_0, 
        m16_2_0, N_5, N_29_i, m37_2_1_1, N_38, N_134_mux, m16_1, m16_2, 
        N_17, N_549, N_125_mux, N_594_1, emflag_cnt_done_0_Z, 
        sig_tapcnt_final_111_3_Z, sig_tapcnt_final_210_3_Z, 
        timeout_fg_3, reset_dly_fg4_4, clkalign_curr_state81_NE_3_Z, 
        N_634_i, N_552_i, N_637, N_653, N_639, N_60, N_523, N_644, 
        N_538_i, N_585_i, no_early_and_late_found_Z, 
        un1_RX_CLK_ALIGN_LOAD5_0_a3_1_1, m122_0_0, tap_cnt9_i_0, 
        un1_early_late_end_set12_3_i_0, m44_0, 
        sig_tapcnt_final_111_4_Z, sig_tapcnt_final_210_4_Z, 
        un1_clkalign_curr_state_1_0_a3_0, emflag_cnt10_i_0, 
        clkalign_curr_state63_NE_3, clkalign_curr_state63_NE_2, 
        clkalign_curr_state63_NE_1, clkalign_curr_state63_NE_0, 
        timeout_fg_4, reset_dly_fg4_6, clkalign_curr_state81_NE_4_Z, 
        N_127_mux, N_619, N_620, N_128_mux, tapcnt_final_0_sqmuxa_1, 
        N_656, N_602_2, N_651, N_657, clkalign_curr_state81, N_27, 
        N_132_mux, N_131_mux, clkalign_curr_state_0_sqmuxa_4_0_a3_0, 
        early_late_start_set5_0_a3_1, emflag_cnt_done_5_Z, 
        un1_early_late_end_set12_1_0_a3_1, emflag_cnt10_i_1, 
        reset_dly_fg4_8, N_490, clkalign_curr_state_1_sqmuxa_1, 
        tapcnt_final_2_sqmuxa_1, N_593, 
        un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0, 
        un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0_0, N_622, N_606_1, 
        N_83, N_138_mux, i22_mux, 
        un1_clkalign_curr_state_1_sqmuxa_5_0_0, 
        un1_clkalign_curr_state_0_sqmuxa_6_0_0_933_1, N_607, N_116, 
        N_93, clkalign_curr_state63, N_143_mux, N_101, 
        emflag_cnt10_i_3, N_118, N_659, N_621, N_594, 
        un1_RX_CLK_ALIGN_LOAD5_0_1, N_3109_mux, N_88, N_25, N_89, 
        N_1835, N_1828, N_1827, N_1249, N_99, N_98, N_97_0, N_96, N_95, 
        N_94, N_93_0, N_92, N_91, N_90, N_89_0, N_88_0, N_87_0, N_86, 
        N_85, N_84, N_83_0, N_82, N_81, N_80, N_79, N_78_0, N_77, N_76, 
        N_75_0, N_74, N_73, N_72, N_71_0, N_70, N_69, N_68, N_67, N_66, 
        N_65, N_64, N_63_0, N_62, N_61_0, N_60_0, N_59, N_58_0, N_57, 
        N_56, N_55_0, N_54, N_53, N_52, N_51, N_50, N_49, N_48, N_47, 
        N_46_0, N_45, N_44, N_43, N_42, N_41, N_40, N_39, N_38_0, N_37, 
        N_36, N_21, N_20, N_19, N_18, N_17_0, N_16, N_15, N_14, N_13, 
        N_12_0;
    
    SLE \cnt[0]  (.D(CO0_0_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(VCC), .ALn(current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND)
        , .LAT(GND), .Q(CO0_0));
    CFG4 #( .INIT(16'hFFBA) )  
        \clkalign_curr_state_ns_5_0_.un1_RX_CLK_ALIGN_LOAD5_0  (.A(
        un1_RX_CLK_ALIGN_LOAD5_0_1), .B(clkalign_curr_state_Z[0]), .C(
        N_606_1), .D(N_607), .Y(un1_RX_CLK_ALIGN_LOAD5_0));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_33 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_63_2_1_co1_15), .S(
        late_found_lsb_63_2_1_wmux_33_S), .Y(
        late_found_lsb_63_2_1_wmux_33_Y), .FCO(
        late_found_lsb_63_2_1_co0_16));
    SLE \late_flags_msb[50]  (.D(late_flags_msb_Z[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[50]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_14 (.A(
        early_found_lsb_126_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[53]), .D(early_flags_lsb_Z[117]), .FCI(
        early_found_lsb_126_2_1_co0_6), .S(
        early_found_lsb_126_2_1_wmux_14_S), .Y(
        early_found_lsb_126_2_1_y3_0), .FCO(
        early_found_lsb_126_2_1_co1_6));
    CFG3 #( .INIT(8'h20) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_2_sqmuxa_1  (.A(
        clkalign_curr_state_d[27]), .B(N_552_i), .C(N_538_i), .Y(
        tapcnt_final_2_sqmuxa_1));
    SLE \late_flags_msb[98]  (.D(late_flags_msb_Z[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[98]));
    CFG4 #( .INIT(16'h8000) )  emflag_cnt_done_5 (.A(emflag_cnt_Z[4]), 
        .B(emflag_cnt_done_0_Z), .C(emflag_cnt_Z[5]), .D(
        emflag_cnt_Z[3]), .Y(emflag_cnt_done_5_Z));
    SLE \early_flags_msb[97]  (.D(early_flags_msb_Z[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[97]));
    CFG3 #( .INIT(8'h80) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0_0  
        (.A(N_627), .B(N_637), .C(N_644), .Y(
        un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0_0));
    SLE \late_flags_lsb[118]  (.D(late_flags_lsb_Z[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[118]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_63_2_1_wmux_43 (.A(
        early_found_lsb_63_2_1_y7_2), .B(early_found_lsb_63_2_1_y5_2), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co1_20), .S(
        early_found_lsb_63_2_1_wmux_43_S), .Y(
        early_found_lsb_63_2_1_y0_19), .FCO(
        early_found_lsb_63_2_1_co0_21));
    CFG2 #( .INIT(4'h2) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_0_sqmuxa_4_0_a3_0  
        (.A(N_656), .B(N_523), .Y(
        clkalign_curr_state_0_sqmuxa_4_0_a3_0));
    SLE \late_flags_msb[14]  (.D(late_flags_msb_Z[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[14]));
    SLE \early_flags_msb[103]  (.D(early_flags_msb_Z[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[103]));
    CFG4 #( .INIT(16'h4A4F) )  \clkalign_curr_state_ns_5_0_.m37_2_1  (
        .A(clkalign_curr_state_Z[1]), .B(N_29_i), .C(m37_2_1_1), .D(
        m37_2_1_1_0), .Y(N_38));
    SLE \late_flags_lsb[124]  (.D(late_flags_lsb_Z[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[124]));
    SLE \late_flags_msb[39]  (.D(late_flags_msb_Z[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[39]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_8 (.A(
        early_found_msb_63_2_1_y0_3), .B(early_found_msb_63_2_1_0_y3), 
        .C(early_found_msb_63_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co0_3), .S(
        early_found_msb_63_2_1_wmux_8_S), .Y(
        early_found_msb_63_2_1_0_y9), .FCO(
        early_found_msb_63_2_1_co1_3));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_38 (.A(
        early_found_lsb_63_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[54]), .D(early_flags_lsb_Z[118]), .FCI(
        early_found_lsb_63_2_1_co0_18), .S(
        early_found_lsb_63_2_1_wmux_38_S), .Y(
        early_found_lsb_63_2_1_y3_2), .FCO(
        early_found_lsb_63_2_1_co1_18));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[14])
        , .D(late_flags_msb_Z[78]), .FCI(late_found_msb_63_2_1_co1_18), 
        .S(late_found_msb_63_2_1_wmux_39_S), .Y(
        late_found_msb_63_2_1_y0_17), .FCO(
        late_found_msb_63_2_1_co0_19));
    SLE \early_flags_lsb[10]  (.D(early_flags_lsb_Z[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[10]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_24 (.A(
        early_found_lsb_63_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[34]), .D(early_flags_lsb_Z[98]), .FCI(
        early_found_lsb_63_2_1_co0_11), .S(
        early_found_lsb_63_2_1_wmux_24_S), .Y(
        early_found_lsb_63_2_1_y1_1), .FCO(
        early_found_lsb_63_2_1_co1_11));
    SLE \early_flags_msb[44]  (.D(early_flags_msb_Z[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[44]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[2]), 
        .D(late_flags_msb_Z[66]), .FCI(late_found_msb_63_2_1_co1_10), 
        .S(late_found_msb_63_2_1_wmux_23_S), .Y(
        late_found_msb_63_2_1_y0_10), .FCO(
        late_found_msb_63_2_1_co0_11));
    SLE \late_flags_lsb[18]  (.D(late_flags_lsb_Z[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[18]));
    SLE \late_flags_msb[26]  (.D(late_flags_msb_Z[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[26]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_20 (.A(
        early_found_lsb_126_2_1_y0_9), .B(early_found_lsb_126_2_1_y3_0)
        , .C(early_found_lsb_126_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_126_2_1_co0_9), .S(
        early_found_lsb_126_2_1_wmux_20_S), .Y(
        early_found_lsb_126_2_1_0_y21), .FCO(
        early_found_lsb_126_2_1_co1_9));
    SLE \early_flags_lsb[49]  (.D(early_flags_lsb_Z[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[49]));
    CFG2 #( .INIT(4'hB) )  
        \clkalign_curr_state_ns_5_0_.un1_RX_CLK_ALIGN_LOAD5_0_o2  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[0]), .Y(
        N_525));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[0]), 
        .D(late_flags_msb_Z[64]), .FCI(VCC), .S(
        late_found_msb_63_2_1_0_wmux_S), .Y(late_found_msb_63_2_1_0_y0)
        , .FCO(late_found_msb_63_2_1_0_co0));
    SLE \late_flags_msb[23]  (.D(late_flags_msb_Z[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[23]));
    CFG3 #( .INIT(8'h27) )  late_found_lsb_127_i (.A(emflag_cnt_Z[0]), 
        .B(N_2094), .C(N_2031), .Y(late_found_lsb_i));
    SLE \late_flags_msb[89]  (.D(late_flags_msb_Z[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[89]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_36 (.A(
        early_found_lsb_63_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[38]), .D(early_flags_lsb_Z[102]), .FCI(
        early_found_lsb_63_2_1_co0_17), .S(
        early_found_lsb_63_2_1_wmux_36_S), .Y(
        early_found_lsb_63_2_1_y1_2), .FCO(
        early_found_lsb_63_2_1_co1_17));
    SLE \late_flags_lsb[123]  (.D(late_flags_lsb_Z[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[123]));
    SLE \early_flags_lsb[50]  (.D(early_flags_lsb_Z[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[50]));
    CFG2 #( .INIT(4'h1) )  sig_tapcnt_final_210_3 (.A(
        early_late_nxt_val_Z[0]), .B(early_late_nxt_val_Z[5]), .Y(
        sig_tapcnt_final_210_3_Z));
    CFG2 #( .INIT(4'h2) )  \clkalign_curr_state_ns_5_0_.m105  (.A(
        N_105), .B(clkalign_curr_state_Z[5]), .Y(
        clkalign_curr_state_ns[3]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_63_2_1_wmux_43 (.A(
        late_found_lsb_63_2_1_y7_2), .B(late_found_lsb_63_2_1_y5_2), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co1_20), .S(
        late_found_lsb_63_2_1_wmux_43_S), .Y(
        late_found_lsb_63_2_1_y0_19), .FCO(
        late_found_lsb_63_2_1_co0_21));
    SLE \early_flags_msb[41]  (.D(early_flags_msb_Z[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[41]));
    SLE \early_flags_msb[52]  (.D(early_flags_msb_Z[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[52]));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_2 (.A(
        early_late_init_val_Z[2]), .B(early_late_nxt_val_Z[2]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_1_Z), .S(
        un2_sig_tapcnt_final_2_cry_2_S), .Y(
        un2_sig_tapcnt_final_2_cry_2_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_2_Z));
    SLE \late_flags_msb[108]  (.D(late_flags_msb_Z[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[108]));
    SLE \early_flags_msb[2]  (.D(early_flags_msb_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[2]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_40 (.A(
        late_found_msb_126_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[47]), .D(late_flags_msb_Z[111]), .FCI(
        late_found_msb_126_2_1_co0_19), .S(
        late_found_msb_126_2_1_wmux_40_S), .Y(
        late_found_msb_126_2_1_y5_2), .FCO(
        late_found_msb_126_2_1_co1_19));
    SLE \early_flags_lsb[65]  (.D(early_flags_lsb_Z[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[65]));
    CFG4 #( .INIT(16'h1000) )  sig_tapcnt_final_210 (.A(
        early_late_nxt_val_Z[2]), .B(early_late_nxt_val_Z[3]), .C(
        sig_tapcnt_final_210_4_Z), .D(sig_tapcnt_final_210_3_Z), .Y(
        sig_tapcnt_final_210_Z));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_cry[4]  (.A(VCC), .B(
        timeout_cnt_Z[4]), .C(GND), .D(GND), .FCI(timeout_cnt_cry_Z[3])
        , .S(timeout_cnt_s[4]), .Y(timeout_cnt_cry_Y[4]), .FCO(
        timeout_cnt_cry_Z[4]));
    SLE \late_flags_lsb[51]  (.D(late_flags_lsb_Z[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[51]));
    SLE \early_flags_msb[46]  (.D(early_flags_msb_Z[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[46]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[22]), .D(early_flags_lsb_Z[86]), .FCI(
        early_found_lsb_63_2_1_co1_17), .S(
        early_found_lsb_63_2_1_wmux_37_S), .Y(
        early_found_lsb_63_2_1_y0_16), .FCO(
        early_found_lsb_63_2_1_co0_18));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_14 (.A(
        early_found_lsb_63_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[52]), .D(early_flags_lsb_Z[116]), .FCI(
        early_found_lsb_63_2_1_co0_6), .S(
        early_found_lsb_63_2_1_wmux_14_S), .Y(
        early_found_lsb_63_2_1_y3_0), .FCO(
        early_found_lsb_63_2_1_co1_6));
    CFG4 #( .INIT(16'hFF59) )  
        \clkalign_curr_state_ns_5_0_.emflag_cnt10_i_1  (.A(
        clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[2]), .C(
        clkalign_curr_state_Z[1]), .D(N_2979), .Y(emflag_cnt10_i_1));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[29])
        , .D(late_flags_lsb_Z[93]), .FCI(late_found_lsb_126_2_1_co1_7), 
        .S(late_found_lsb_126_2_1_wmux_17_S), .Y(
        late_found_lsb_126_2_1_y0_8), .FCO(
        late_found_lsb_126_2_1_co0_8));
    SLE \late_flags_msb[106]  (.D(late_flags_msb_Z[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[106]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[1])
        , .D(early_flags_msb_Z[65]), .FCI(VCC), .S(
        early_found_msb_126_2_1_0_wmux_S), .Y(
        early_found_msb_126_2_1_0_y0), .FCO(
        early_found_msb_126_2_1_0_co0));
    SLE \early_flags_msb[7]  (.D(early_flags_msb_Z[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[7]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[25])
        , .D(late_flags_msb_Z[89]), .FCI(late_found_msb_126_2_1_co1_1), 
        .S(late_found_msb_126_2_1_wmux_5_S), .Y(
        late_found_msb_126_2_1_y0_2), .FCO(
        late_found_msb_126_2_1_co0_2));
    SLE \early_flags_msb[94]  (.D(early_flags_msb_Z[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[94]));
    SLE \early_flags_lsb[25]  (.D(early_flags_lsb_Z[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[25]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_12 (.A(
        late_found_lsb_126_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[37]), .D(late_flags_lsb_Z[101]), .FCI(
        late_found_lsb_126_2_1_co0_5), .S(
        late_found_lsb_126_2_1_wmux_12_S), .Y(
        late_found_lsb_126_2_1_y1_0), .FCO(
        late_found_lsb_126_2_1_co1_5));
    SLE \late_flags_lsb[55]  (.D(late_flags_lsb_Z[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[55]));
    SLE \early_flags_msb[111]  (.D(early_flags_msb_Z[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[111]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_22 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_63_2_1_co0_10), .S(
        early_found_msb_63_2_1_wmux_22_S), .Y(
        early_found_msb_63_2_1_wmux_22_Y), .FCO(
        early_found_msb_63_2_1_co1_10));
    SLE \timeout_cnt[7]  (.D(timeout_cnt_s_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[7]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_32 (.A(
        early_found_msb_126_2_1_y0_14), .B(
        early_found_msb_126_2_1_y3_1), .C(early_found_msb_126_2_1_y1_1)
        , .D(emflag_cnt_Z[3]), .FCI(early_found_msb_126_2_1_co0_15), 
        .S(early_found_msb_126_2_1_wmux_32_S), .Y(
        early_found_msb_126_2_1_0_y33), .FCO(
        early_found_msb_126_2_1_co1_15));
    SLE \late_flags_lsb[114]  (.D(late_flags_lsb_Z[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[114]));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNIUBO91[0]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[0]), 
        .D(GND), .FCI(tapcnt_offset_cry_cy), .S(tapcnt_offset_s[0]), 
        .Y(tapcnt_offset_RNIUBO91_Y[0]), .FCO(tapcnt_offset_cry[0]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_20 (.A(
        late_found_msb_126_2_1_y0_9), .B(late_found_msb_126_2_1_y3_0), 
        .C(late_found_msb_126_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co0_9), .S(
        late_found_msb_126_2_1_wmux_20_S), .Y(
        late_found_msb_126_2_1_0_y21), .FCO(
        late_found_msb_126_2_1_co1_9));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[25]), .D(early_flags_msb_Z[89]), .FCI(
        early_found_msb_126_2_1_co1_1), .S(
        early_found_msb_126_2_1_wmux_5_S), .Y(
        early_found_msb_126_2_1_y0_2), .FCO(
        early_found_msb_126_2_1_co0_2));
    CFG4 #( .INIT(16'h3A30) )  \clkalign_curr_state_ns_5_0_.m86_1  (.A(
        calc_done_Z), .B(clkalign_curr_state_Z[0]), .C(
        clkalign_curr_state_Z[1]), .D(N_19_i), .Y(m86_1_0));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_12 (.A(
        early_found_msb_63_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[36]), .D(early_flags_msb_Z[100]), .FCI(
        early_found_msb_63_2_1_co0_5), .S(
        early_found_msb_63_2_1_wmux_12_S), .Y(
        early_found_msb_63_2_1_y1_0), .FCO(
        early_found_msb_63_2_1_co1_5));
    SLE \early_flags_msb[48]  (.D(early_flags_msb_Z[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[48]));
    SLE \late_flags_msb[77]  (.D(late_flags_msb_Z[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[77]));
    SLE \late_flags_msb[99]  (.D(late_flags_msb_Z[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[99]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[17]), .D(early_flags_msb_Z[81]), .FCI(
        early_found_msb_126_2_1_0_co1), .S(
        early_found_msb_126_2_1_wmux_1_S), .Y(
        early_found_msb_126_2_1_y0_0), .FCO(
        early_found_msb_126_2_1_co0_0));
    SLE \late_flags_lsb[20]  (.D(late_flags_lsb_Z[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[20]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_33 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_126_2_1_co1_15), .S(
        late_found_msb_126_2_1_wmux_33_S), .Y(
        late_found_msb_126_2_1_wmux_33_Y), .FCO(
        late_found_msb_126_2_1_co0_16));
    SLE \early_flags_msb[91]  (.D(early_flags_msb_Z[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[91]));
    SLE \early_flags_lsb[118]  (.D(early_flags_lsb_Z[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[118]));
    ARI1 #( .INIT(20'h0F588) )  
        \clkalign_curr_state_ns_5_0_.m70_1_0_wmux_0  (.A(m70_1_0_y0), 
        .B(clkalign_curr_state_Z[3]), .C(N_63), .D(i18_mux), .FCI(
        m70_1_0_co0), .S(m70_1_0_wmux_0_S), .Y(N_71), .FCO(m70_1_0_co1)
        );
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[15])
        , .D(late_flags_msb_Z[79]), .FCI(late_found_msb_126_2_1_co1_18)
        , .S(late_found_msb_126_2_1_wmux_39_S), .Y(
        late_found_msb_126_2_1_y0_17), .FCO(
        late_found_msb_126_2_1_co0_19));
    SLE \early_late_end_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[5]));
    SLE no_early_and_late_found_msb_d (.D(
        no_early_and_late_found_msb_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(no_early_and_late_found_msb_d_Z));
    CFG2 #( .INIT(4'h1) )  
        \clkalign_curr_state_ns_5_0_.early_late_init_set5_0_a2  (.A(
        clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[2]), .Y(
        N_637));
    SLE \late_flags_lsb[113]  (.D(late_flags_lsb_Z[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[113]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_1 
        (.A(early_late_nxt_val_Z[1]), .B(early_late_init_val_Z[1]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_0_Z), 
        .S(early_late_init_nxt_val_status5_cry_1_S), .Y(
        early_late_init_nxt_val_status5_cry_1_Y), .FCO(
        early_late_init_nxt_val_status5_cry_1_Z));
    SLE \early_flags_lsb[87]  (.D(early_flags_lsb_Z[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[87]));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_0 (.A(
        early_late_end_val_Z[0]), .B(early_late_start_val_Z[0]), .C(
        GND), .D(GND), .FCI(GND), .S(un3_sig_tapcnt_final_1_cry_0_S), 
        .Y(un3_sig_tapcnt_final_1_cry_0_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_0_Z));
    SLE \early_flags_msb[96]  (.D(early_flags_msb_Z[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[96]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_63_2_1_wmux_7 (.A(
        early_found_lsb_63_2_1_0_y7), .B(early_found_lsb_63_2_1_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co1_2), .S(
        early_found_lsb_63_2_1_wmux_7_S), .Y(
        early_found_lsb_63_2_1_y0_3), .FCO(
        early_found_lsb_63_2_1_co0_3));
    SLE \late_flags_lsb[80]  (.D(late_flags_lsb_Z[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[80]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[6]  (.A(
        tapcnt_final_11_iv_1[6]), .B(tapcnt_final_11_iv_0[6]), .Y(
        tapcnt_final_11[6]));
    CFG3 #( .INIT(8'h2F) )  \clkalign_curr_state_ns_5_0_.m67  (.A(N_61)
        , .B(no_early_and_late_found_Z), .C(clkalign_curr_state_Z[1]), 
        .Y(N_138_mux));
    CFG2 #( .INIT(4'h9) )  \clkalign_curr_state_ns_5_0_.m16_1  (.A(
        clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[1]), .Y(
        m16_1));
    SLE \late_flags_lsb[19]  (.D(late_flags_lsb_Z[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[19]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.RX_CLK_ALIGN_DONE5  (.A(
        timeout_fg), .B(clk_align_done_Z), .Y(RX_CLK_ALIGN_DONE5));
    SLE \late_flags_lsb[48]  (.D(late_flags_lsb_Z[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[48]));
    SLE \early_flags_lsb[125]  (.D(early_flags_lsb_Z[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[125]));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[1]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[1]), .D(GND), .FCI(
        tap_cnt_cry_Z[0]), .S(tap_cnt_s[1]), .Y(tap_cnt_cry_Y[1]), 
        .FCO(tap_cnt_cry_Z[1]));
    CFG4 #( .INIT(16'hC0EA) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_8_0_o2  
        (.A(N_627), .B(clkalign_curr_state_Z[4]), .C(N_656), .D(N_523), 
        .Y(N_526));
    SLE early_or_late_found_lsb_d (.D(early_or_late_found_lsb_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_or_late_found_lsb_d_Z));
    SLE \early_late_end_val[7]  (.D(emflag_cnt_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[7]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_16 (.A(
        late_found_lsb_63_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[44]), .D(late_flags_lsb_Z[108]), .FCI(
        late_found_lsb_63_2_1_co0_7), .S(
        late_found_lsb_63_2_1_wmux_16_S), .Y(
        late_found_lsb_63_2_1_y5_0), .FCO(late_found_lsb_63_2_1_co1_7));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[4]), 
        .D(late_flags_msb_Z[68]), .FCI(late_found_msb_63_2_1_co1_4), 
        .S(late_found_msb_63_2_1_wmux_11_S), .Y(
        late_found_msb_63_2_1_y0_5), .FCO(late_found_msb_63_2_1_co0_5));
    SLE \late_flags_msb[74]  (.D(late_flags_msb_Z[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[74]));
    SLE \early_flags_msb[55]  (.D(early_flags_msb_Z[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[55]));
    CFG3 #( .INIT(8'h80) )  \clkalign_curr_state_ns_5_0_.m81  (.A(
        clkalign_curr_state_Z[4]), .B(emflag_cnt_done_d_Z), .C(
        clkalign_curr_state_Z[0]), .Y(N_82_i));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_63_2_1_wmux_31 (.A(
        late_found_lsb_63_2_1_y7_1), .B(late_found_lsb_63_2_1_y5_1), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co1_14), .S(
        late_found_lsb_63_2_1_wmux_31_S), .Y(
        late_found_lsb_63_2_1_y0_14), .FCO(
        late_found_lsb_63_2_1_co0_15));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[21]), .D(early_flags_lsb_Z[85]), .FCI(
        early_found_lsb_126_2_1_co1_5), .S(
        early_found_lsb_126_2_1_wmux_13_S), .Y(
        early_found_lsb_126_2_1_y0_6), .FCO(
        early_found_lsb_126_2_1_co0_6));
    SLE \clkalign_curr_state[1]  (.D(clkalign_curr_state_ns[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(clkalign_curr_state_Z[1]));
    SLE \timeout_cnt[4]  (.D(timeout_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[4]));
    SLE \late_flags_msb[60]  (.D(late_flags_msb_Z[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[60]));
    SLE \early_flags_msb[98]  (.D(early_flags_msb_Z[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[98]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_4 (.A(
        late_found_lsb_126_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[41]), .D(late_flags_lsb_Z[105]), .FCI(
        late_found_lsb_126_2_1_co0_1), .S(
        late_found_lsb_126_2_1_wmux_4_S), .Y(
        late_found_lsb_126_2_1_0_y5), .FCO(
        late_found_lsb_126_2_1_co1_1));
    SLE \late_flags_lsb[120]  (.D(late_flags_lsb_Z[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[120]));
    SLE \wait_cnt[2]  (.D(wait_cnt_3[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(wait_cnt_Z[2]));
    SLE \early_late_end_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[2]));
    SLE \tap_cnt[7]  (.D(tap_cnt_s_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[7]));
    SLE \early_flags_msb[119]  (.D(early_flags_msb_Z[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[119]));
    SLE \late_flags_msb[122]  (.D(late_flags_msb_Z[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[122]));
    SLE \late_flags_lsb[76]  (.D(late_flags_lsb_Z[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[76]));
    CFG2 #( .INIT(4'h8) )  \clkalign_curr_state_ns_5_0_.m2_e  (.A(
        CO0_0), .B(cnt_Z[1]), .Y(N_125_mux));
    SLE \late_flags_lsb[73]  (.D(late_flags_lsb_Z[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[73]));
    SLE \early_flags_msb[79]  (.D(early_flags_msb_Z[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[79]));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_2 (.A(
        early_late_end_val_Z[2]), .B(early_late_start_val_Z[2]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_1_Z), .S(
        un3_sig_tapcnt_final_1_cry_2_S), .Y(
        un3_sig_tapcnt_final_1_cry_2_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_2_Z));
    SLE \early_flags_msb[10]  (.D(early_flags_msb_Z[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[10]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_36 (.A(
        late_found_lsb_126_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[39]), .D(late_flags_lsb_Z[103]), .FCI(
        late_found_lsb_126_2_1_co0_17), .S(
        late_found_lsb_126_2_1_wmux_36_S), .Y(
        late_found_lsb_126_2_1_y1_2), .FCO(
        late_found_lsb_126_2_1_co1_17));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_18 (.A(
        early_found_msb_126_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[61]), .D(early_flags_msb_Z[125]), .FCI(
        early_found_msb_126_2_1_co0_8), .S(
        early_found_msb_126_2_1_wmux_18_S), .Y(
        early_found_msb_126_2_1_y7_0), .FCO(
        early_found_msb_126_2_1_co1_8));
    SLE \late_flags_lsb[119]  (.D(late_flags_lsb_Z[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[119]));
    SLE \early_flags_lsb[112]  (.D(early_flags_lsb_Z[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[112]));
    SLE \early_flags_lsb[105]  (.D(early_flags_lsb_Z[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[105]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[0]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[0]), .D(early_late_start_val_Z[0]), 
        .Y(tapcnt_final_11_iv_0[0]));
    CFG4 #( .INIT(16'h4000) )  
        \clkalign_curr_state_ns_5_0_.RX_CLK_ALIGN_LOAD5_0_a3_0_1  (.A(
        N_549), .B(N_2979), .C(N_125_mux), .D(calc_done_Z), .Y(N_594_1)
        );
    CFG3 #( .INIT(8'hF2) )  \clkalign_curr_state_ns_5_0_.m86  (.A(
        m86_1_0), .B(clkalign_curr_state_Z[4]), .C(m86_2), .Y(N_87));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[6]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_7_S), 
        .Y(sig_tapcnt_final_1_3_Z[6]));
    SLE \early_flags_lsb[0]  (.D(early_flags_lsb_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[0]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_32 (.A(
        early_found_lsb_126_2_1_y0_14), .B(
        early_found_lsb_126_2_1_y3_1), .C(early_found_lsb_126_2_1_y1_1)
        , .D(emflag_cnt_Z[3]), .FCI(early_found_lsb_126_2_1_co0_15), 
        .S(early_found_lsb_126_2_1_wmux_32_S), .Y(
        early_found_lsb_126_2_1_0_y33), .FCO(
        early_found_lsb_126_2_1_co1_15));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[5])
        , .D(early_flags_lsb_Z[69]), .FCI(
        early_found_lsb_126_2_1_co1_4), .S(
        early_found_lsb_126_2_1_wmux_11_S), .Y(
        early_found_lsb_126_2_1_y0_5), .FCO(
        early_found_lsb_126_2_1_co0_5));
    SLE \late_flags_lsb[38]  (.D(late_flags_lsb_Z[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[38]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_63_2_1_wmux_43 (.A(
        early_found_msb_63_2_1_y7_2), .B(early_found_msb_63_2_1_y5_2), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co1_20), .S(
        early_found_msb_63_2_1_wmux_43_S), .Y(
        early_found_msb_63_2_1_y0_19), .FCO(
        early_found_msb_63_2_1_co0_21));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_21 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_63_2_1_co1_9), .S(
        late_found_msb_63_2_1_wmux_21_S), .Y(
        late_found_msb_63_2_1_wmux_21_Y), .FCO(
        late_found_msb_63_2_1_co0_10));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_6 (.A(
        late_found_msb_63_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[56]), .D(late_flags_msb_Z[120]), .FCI(
        late_found_msb_63_2_1_co0_2), .S(
        late_found_msb_63_2_1_wmux_6_S), .Y(late_found_msb_63_2_1_0_y7)
        , .FCO(late_found_msb_63_2_1_co1_2));
    SLE \early_flags_msb[33]  (.D(early_flags_msb_Z[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[33]));
    SLE RX_CLK_ALIGN_CLR_FLGS (.D(N_2939), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_0_sqmuxa_8_0), .ALn(current_state_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_34 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_126_2_1_co0_16), .S(
        late_found_lsb_126_2_1_wmux_34_S), .Y(
        late_found_lsb_126_2_1_wmux_34_Y), .FCO(
        late_found_lsb_126_2_1_co1_16));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[13]), .D(early_flags_lsb_Z[77]), .FCI(
        early_found_lsb_126_2_1_co1_6), .S(
        early_found_lsb_126_2_1_wmux_15_S), .Y(
        early_found_lsb_126_2_1_y0_7), .FCO(
        early_found_lsb_126_2_1_co0_7));
    SLE \early_flags_lsb[84]  (.D(early_flags_lsb_Z[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[84]));
    CFG3 #( .INIT(8'hD8) )  \clkalign_curr_state_ns_5_0_.m68  (.A(
        clkalign_curr_state_Z[4]), .B(N_138_mux), .C(i22_mux), .Y(
        i18_mux));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_28 (.A(
        early_found_msb_63_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[42]), .D(early_flags_msb_Z[106]), .FCI(
        early_found_msb_63_2_1_co0_13), .S(
        early_found_msb_63_2_1_wmux_28_S), .Y(
        early_found_msb_63_2_1_y5_1), .FCO(
        early_found_msb_63_2_1_co1_13));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNI4TBR4[5]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[5]), 
        .D(GND), .FCI(tapcnt_offset_cry[4]), .S(tapcnt_offset_s[5]), 
        .Y(tapcnt_offset_RNI4TBR4_Y[5]), .FCO(tapcnt_offset_cry[5]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_2 (.A(
        late_found_lsb_126_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[49]), .D(late_flags_lsb_Z[113]), .FCI(
        late_found_lsb_126_2_1_co0_0), .S(
        late_found_lsb_126_2_1_wmux_2_S), .Y(
        late_found_lsb_126_2_1_0_y3), .FCO(
        late_found_lsb_126_2_1_co1_0));
    SLE \early_flags_lsb[119]  (.D(early_flags_lsb_Z[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[119]));
    SLE \late_flags_msb[11]  (.D(late_flags_msb_Z[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[11]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_18 (.A(
        early_found_msb_63_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[60]), .D(early_flags_msb_Z[124]), .FCI(
        early_found_msb_63_2_1_co0_8), .S(
        early_found_msb_63_2_1_wmux_18_S), .Y(
        early_found_msb_63_2_1_y7_0), .FCO(
        early_found_msb_63_2_1_co1_8));
    CFG4 #( .INIT(16'h8000) )  
        \clkalign_curr_state_ns_5_0_.reset_dly_fg4  (.A(rst_cnt_Z[0]), 
        .B(reset_dly_fg4_8), .C(rst_cnt_Z[1]), .D(reset_dly_fg4_4), .Y(
        reset_dly_fg4));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[30])
        , .D(late_flags_lsb_Z[94]), .FCI(late_found_lsb_63_2_1_co1_19), 
        .S(late_found_lsb_63_2_1_wmux_41_S), .Y(
        late_found_lsb_63_2_1_y0_18), .FCO(
        late_found_lsb_63_2_1_co0_20));
    CFG3 #( .INIT(8'h40) )  
        \clkalign_curr_state_ns_5_0_.un1_RX_CLK_ALIGN_LOAD5_0_a3_0_1  
        (.A(N_523), .B(N_642), .C(N_627), .Y(N_606_1));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_32 (.A(
        early_found_msb_63_2_1_y0_14), .B(early_found_msb_63_2_1_y3_1), 
        .C(early_found_msb_63_2_1_y1_1), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co0_15), .S(
        early_found_msb_63_2_1_wmux_32_S), .Y(
        early_found_msb_63_2_1_0_y33), .FCO(
        early_found_msb_63_2_1_co1_15));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[18]), .D(early_flags_lsb_Z[82]), .FCI(
        early_found_lsb_63_2_1_co1_11), .S(
        early_found_lsb_63_2_1_wmux_25_S), .Y(
        early_found_lsb_63_2_1_y0_11), .FCO(
        early_found_lsb_63_2_1_co0_12));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_26 (.A(
        early_found_msb_63_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[50]), .D(early_flags_msb_Z[114]), .FCI(
        early_found_msb_63_2_1_co0_12), .S(
        early_found_msb_63_2_1_wmux_26_S), .Y(
        early_found_msb_63_2_1_y3_1), .FCO(
        early_found_msb_63_2_1_co1_12));
    CLKINT RX_CLK_ALIGN_DONE_rep_RNIOGJF (.A(RX_CLK_ALIGN_DONE_rep_Z), 
        .Y(RX_CLK_ALIGN_DONE_arst));
    CFG4 #( .INIT(16'hF020) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_i_0[0]  (.A(N_659), .B(
        clkalign_curr_state_Z[0]), .C(wait_cnt_Z[0]), .D(
        wait_cnt_3_i_a3_2_0[0]), .Y(wait_cnt_3_i_0[0]));
    ARI1 #( .INIT(20'h0CEC2) )  late_found_msb_126_2_1_wmux_10 (.A(
        late_found_msb_126_2_1_0_y21), .B(late_found_msb_126_2_1_0_y9), 
        .C(emflag_cnt_Z[2]), .D(emflag_cnt_Z[1]), .FCI(
        late_found_msb_126_2_1_co0_4), .S(
        late_found_msb_126_2_1_wmux_10_S), .Y(
        late_found_msb_126_2_1_y0_4), .FCO(
        late_found_msb_126_2_1_co1_4));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_26 (.A(
        early_found_msb_126_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[51]), .D(early_flags_msb_Z[115]), .FCI(
        early_found_msb_126_2_1_co0_12), .S(
        early_found_msb_126_2_1_wmux_26_S), .Y(
        early_found_msb_126_2_1_y3_1), .FCO(
        early_found_msb_126_2_1_co1_12));
    SLE \early_flags_lsb[9]  (.D(early_flags_lsb_Z[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[9]));
    SLE \early_flags_lsb[81]  (.D(early_flags_lsb_Z[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[81]));
    CFG4 #( .INIT(16'h0001) )  sig_tapcnt_final_111_4 (.A(
        early_late_end_val_Z[7]), .B(early_late_end_val_Z[6]), .C(
        early_late_end_val_Z[5]), .D(early_late_end_val_Z[4]), .Y(
        sig_tapcnt_final_111_4_Z));
    ARI1 #( .INIT(20'h0CEC2) )  early_found_msb_126_2_1_wmux_10 (.A(
        early_found_msb_126_2_1_0_y21), .B(
        early_found_msb_126_2_1_0_y9), .C(emflag_cnt_Z[2]), .D(
        emflag_cnt_Z[1]), .FCI(early_found_msb_126_2_1_co0_4), .S(
        early_found_msb_126_2_1_wmux_10_S), .Y(
        early_found_msb_126_2_1_y0_4), .FCO(
        early_found_msb_126_2_1_co1_4));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_16 (.A(
        early_found_msb_63_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[44]), .D(early_flags_msb_Z[108]), .FCI(
        early_found_msb_63_2_1_co0_7), .S(
        early_found_msb_63_2_1_wmux_16_S), .Y(
        early_found_msb_63_2_1_y5_0), .FCO(
        early_found_msb_63_2_1_co1_7));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_8 (.A(
        early_found_lsb_63_2_1_y0_3), .B(early_found_lsb_63_2_1_0_y3), 
        .C(early_found_lsb_63_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co0_3), .S(
        early_found_lsb_63_2_1_wmux_8_S), .Y(
        early_found_lsb_63_2_1_0_y9), .FCO(
        early_found_lsb_63_2_1_co1_3));
    SLE \late_flags_msb[15]  (.D(late_flags_msb_Z[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[15]));
    CFG3 #( .INIT(8'h20) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_1_sqmuxa_1_0_a3  
        (.A(N_602_2), .B(PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), .C(
        N_2979), .Y(clkalign_curr_state_1_sqmuxa_1));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_126_2_1_wmux_7 (.A(
        early_found_msb_126_2_1_0_y7), .B(early_found_msb_126_2_1_0_y5)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_126_2_1_co1_2), .S(
        early_found_msb_126_2_1_wmux_7_S), .Y(
        early_found_msb_126_2_1_y0_3), .FCO(
        early_found_msb_126_2_1_co0_3));
    SLE \early_flags_lsb[86]  (.D(early_flags_lsb_Z[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[86]));
    SLE \timeout_cnt[3]  (.D(timeout_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[3]));
    CFG2 #( .INIT(4'h2) )  \clkalign_curr_state_ns_5_0_.m59  (.A(
        clkalign_curr_state_Z[0]), .B(emflag_cnt_done_d_Z), .Y(N_60));
    SLE \late_flags_lsb[110]  (.D(late_flags_lsb_Z[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[110]));
    SLE \early_flags_lsb[40]  (.D(early_flags_lsb_Z[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[40]));
    SLE \late_flags_lsb[49]  (.D(late_flags_lsb_Z[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[49]));
    SLE \late_flags_msb[112]  (.D(late_flags_msb_Z[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[112]));
    SLE \late_flags_msb[0]  (.D(late_flags_msb_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[0]));
    SLE \timeout_cnt[1]  (.D(timeout_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[1]));
    SLE \late_flags_msb[20]  (.D(late_flags_msb_Z[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[20]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[10]), .D(early_flags_msb_Z[74]), .FCI(
        early_found_msb_63_2_1_co1_12), .S(
        early_found_msb_63_2_1_wmux_27_S), .Y(
        early_found_msb_63_2_1_y0_12), .FCO(
        early_found_msb_63_2_1_co0_13));
    SLE \late_flags_msb[109]  (.D(late_flags_msb_Z[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[109]));
    CFG4 #( .INIT(16'h7DBE) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state63_NE_3  (.A(
        tapcnt_final_Z[0]), .B(tapcnt_final_Z[7]), .C(tap_cnt_Z[7]), 
        .D(tap_cnt_Z[0]), .Y(clkalign_curr_state63_NE_3));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[3]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[3]), .D(GND), .FCI(
        emflag_cnt_cry_Z[2]), .S(emflag_cnt_s[3]), .Y(
        emflag_cnt_cry_Y[3]), .FCO(emflag_cnt_cry_Z[3]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[28]), .D(early_flags_msb_Z[92]), .FCI(
        early_found_msb_63_2_1_co1_7), .S(
        early_found_msb_63_2_1_wmux_17_S), .Y(
        early_found_msb_63_2_1_y0_8), .FCO(
        early_found_msb_63_2_1_co0_8));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[30]), .D(early_flags_lsb_Z[94]), .FCI(
        early_found_lsb_63_2_1_co1_19), .S(
        early_found_lsb_63_2_1_wmux_41_S), .Y(
        early_found_lsb_63_2_1_y0_18), .FCO(
        early_found_lsb_63_2_1_co0_20));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[12]), .D(early_flags_lsb_Z[76]), .FCI(
        early_found_lsb_63_2_1_co1_6), .S(
        early_found_lsb_63_2_1_wmux_15_S), .Y(
        early_found_lsb_63_2_1_y0_7), .FCO(
        early_found_lsb_63_2_1_co0_7));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[4]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[4]), .D(early_late_start_val_Z[4]), 
        .Y(tapcnt_final_11_iv_0[4]));
    SLE \early_flags_lsb[7]  (.D(early_flags_lsb_Z[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[7]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_33 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_126_2_1_co1_15), .S(
        early_found_msb_126_2_1_wmux_33_S), .Y(
        early_found_msb_126_2_1_wmux_33_Y), .FCO(
        early_found_msb_126_2_1_co0_16));
    SLE \late_flags_msb[58]  (.D(late_flags_msb_Z[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[58]));
    SLE \early_flags_msb[42]  (.D(early_flags_msb_Z[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[42]));
    CFG4 #( .INIT(16'h4000) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_11_0_a3  
        (.A(N_525), .B(start_trng_fg_Z), .C(N_627), .D(N_637), .Y(
        N_585_i));
    SLE \early_flags_lsb[114]  (.D(early_flags_lsb_Z[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[114]));
    SLE early_found_msb_d (.D(early_found_msb), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_found_msb_d_Z));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[2]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[2]), .D(early_late_start_val_Z[2]), 
        .Y(tapcnt_final_11_iv_0[2]));
    SLE \early_flags_lsb[88]  (.D(early_flags_lsb_Z[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[88]));
    CFG3 #( .INIT(8'hB8) )  \clkalign_curr_state_ns_5_0_.m16_2_1  (.A(
        m16_2_0), .B(clkalign_curr_state_Z[2]), .C(m16_2), .Y(N_17));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_63_2_1_wmux_19 (.A(
        late_found_lsb_63_2_1_y7_0), .B(late_found_lsb_63_2_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co1_8), .S(
        late_found_lsb_63_2_1_wmux_19_S), .Y(
        late_found_lsb_63_2_1_y0_9), .FCO(late_found_lsb_63_2_1_co0_9));
    CFG3 #( .INIT(8'h13) )  \clkalign_curr_state_ns_5_0_.N_511_i_1  (
        .A(clkalign_curr_state_Z[5]), .B(clkalign_curr_state_Z[3]), .C(
        clkalign_curr_state_Z[0]), .Y(N_511_i_1));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNINF6N2[2]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[2]), 
        .D(GND), .FCI(tapcnt_offset_cry[1]), .S(tapcnt_offset_s[2]), 
        .Y(tapcnt_offset_RNINF6N2_Y[2]), .FCO(tapcnt_offset_cry[2]));
    SLE \late_flags_lsb[8]  (.D(late_flags_lsb_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[8]));
    SLE \late_flags_lsb[39]  (.D(late_flags_lsb_Z[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[39]));
    CFG4 #( .INIT(16'h880A) )  \clkalign_curr_state_ns_5_0_.m28  (.A(
        clkalign_curr_state_Z[4]), .B(N_27), .C(rx_trng_done_Z), .D(
        clkalign_curr_state_Z[0]), .Y(N_29_i));
    SLE \early_flags_msb[63]  (.D(early_flags_msb_Z[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[63]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[1]), 
        .D(late_flags_lsb_Z[65]), .FCI(VCC), .S(
        late_found_lsb_126_2_1_0_wmux_S), .Y(
        late_found_lsb_126_2_1_0_y0), .FCO(
        late_found_lsb_126_2_1_0_co0));
    CFG3 #( .INIT(8'h20) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_end_set12_1_0_a3_1  
        (.A(N_639), .B(N_525), .C(N_627), .Y(
        un1_early_late_end_set12_1_0_a3_1));
    CFG4 #( .INIT(16'hF7FF) )  clkalign_curr_state81_NE_4 (.A(
        tapcnt_offset_Z[4]), .B(tapcnt_offset_Z[3]), .C(
        tapcnt_offset_Z[1]), .D(tapcnt_offset_Z[0]), .Y(
        clkalign_curr_state81_NE_4_Z));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_7 (.A(
        early_late_init_val_Z[7]), .B(early_late_nxt_val_Z[7]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_6_Z), .S(
        un2_sig_tapcnt_final_2_cry_7_S), .Y(
        un2_sig_tapcnt_final_2_cry_7_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_7_Z));
    SLE \early_flags_lsb[17]  (.D(early_flags_lsb_Z[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[17]));
    CFG4 #( .INIT(16'h00BF) )  \clkalign_curr_state_ns_5_0_.m111  (.A(
        early_or_late_found_Z), .B(no_early_and_late_found_Z), .C(N_60)
        , .D(clkalign_curr_state_Z[4]), .Y(N_137_mux));
    CFG3 #( .INIT(8'h7F) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s5_0_a3  (.A(
        N_627), .B(N_644), .C(N_2979), .Y(N_673_i));
    CFG1 #( .INIT(2'h1) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s9_0_a3_RNITJ81  
        (.A(clkalign_curr_state_s9_0_a3), .Y(N_677_i));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_32 (.A(
        late_found_msb_63_2_1_y0_14), .B(late_found_msb_63_2_1_y3_1), 
        .C(late_found_msb_63_2_1_y1_1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co0_15), .S(
        late_found_msb_63_2_1_wmux_32_S), .Y(
        late_found_msb_63_2_1_0_y33), .FCO(
        late_found_msb_63_2_1_co1_15));
    SLE \early_flags_lsb[57]  (.D(early_flags_lsb_Z[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[57]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_38 (.A(
        early_found_msb_63_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[54]), .D(early_flags_msb_Z[118]), .FCI(
        early_found_msb_63_2_1_co0_18), .S(
        early_found_msb_63_2_1_wmux_38_S), .Y(
        early_found_msb_63_2_1_y3_2), .FCO(
        early_found_msb_63_2_1_co1_18));
    VCC VCC_Z (.Y(VCC));
    SLE early_late_start_set (.D(clkalign_curr_state_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(early_late_start_set_Z));
    CFG4 #( .INIT(16'h7BDE) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state63_NE_1  (.A(
        tapcnt_final_Z[4]), .B(tapcnt_final_Z[3]), .C(tap_cnt_Z[4]), 
        .D(tap_cnt_Z[3]), .Y(clkalign_curr_state63_NE_1));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[17])
        , .D(late_flags_lsb_Z[81]), .FCI(late_found_lsb_126_2_1_0_co1), 
        .S(late_found_lsb_126_2_1_wmux_1_S), .Y(
        late_found_lsb_126_2_1_y0_0), .FCO(
        late_found_lsb_126_2_1_co0_0));
    SLE \early_late_start_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[3]));
    CFG3 #( .INIT(8'h40) )  
        \clkalign_curr_state_ns_5_0_.early_late_init_set5_0_a3_0  (.A(
        N_533), .B(N_637), .C(N_644), .Y(N_593));
    SLE \early_flags_msb[92]  (.D(early_flags_msb_Z[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[92]));
    SLE \early_late_start_val[7]  (.D(emflag_cnt_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[7]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[19]), .D(early_flags_msb_Z[83]), .FCI(
        early_found_msb_126_2_1_co1_11), .S(
        early_found_msb_126_2_1_wmux_25_S), .Y(
        early_found_msb_126_2_1_y0_11), .FCO(
        early_found_msb_126_2_1_co0_12));
    SLE \tapcnt_offset[0]  (.D(tapcnt_offset_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[0]));
    ARI1 #( .INIT(20'h0EA4A) )  late_found_msb_126_2_1_wmux_9 (.A(
        late_found_msb_126_2_1_0_y45), .B(late_found_msb_126_2_1_y0_4), 
        .C(late_found_msb_126_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        late_found_msb_126_2_1_co1_3), .S(
        late_found_msb_126_2_1_wmux_9_S), .Y(N_2348), .FCO(
        late_found_msb_126_2_1_co0_4));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_36 (.A(
        early_found_msb_63_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[38]), .D(early_flags_msb_Z[102]), .FCI(
        early_found_msb_63_2_1_co0_17), .S(
        early_found_msb_63_2_1_wmux_36_S), .Y(
        early_found_msb_63_2_1_y1_2), .FCO(
        early_found_msb_63_2_1_co1_17));
    SLE \tap_cnt[6]  (.D(tap_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[6]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_26 (.A(
        late_found_lsb_63_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[50]), .D(late_flags_lsb_Z[114]), .FCI(
        late_found_lsb_63_2_1_co0_12), .S(
        late_found_lsb_63_2_1_wmux_26_S), .Y(
        late_found_lsb_63_2_1_y3_1), .FCO(late_found_lsb_63_2_1_co1_12)
        );
    SLE \late_flags_msb[71]  (.D(late_flags_msb_Z[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[71]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[11]), .D(early_flags_lsb_Z[75]), .FCI(
        early_found_lsb_126_2_1_co1_12), .S(
        early_found_lsb_126_2_1_wmux_27_S), .Y(
        early_found_lsb_126_2_1_y0_12), .FCO(
        early_found_lsb_126_2_1_co0_13));
    ARI1 #( .INIT(20'h0EA4A) )  early_found_lsb_63_2_1_wmux_9 (.A(
        early_found_lsb_63_2_1_0_y45), .B(early_found_lsb_63_2_1_y0_4), 
        .C(early_found_lsb_63_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        early_found_lsb_63_2_1_co1_3), .S(
        early_found_lsb_63_2_1_wmux_9_S), .Y(N_1904), .FCO(
        early_found_lsb_63_2_1_co0_4));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[24])
        , .D(late_flags_lsb_Z[88]), .FCI(late_found_lsb_63_2_1_co1_1), 
        .S(late_found_lsb_63_2_1_wmux_5_S), .Y(
        late_found_lsb_63_2_1_y0_2), .FCO(late_found_lsb_63_2_1_co0_2));
    CFG2 #( .INIT(4'h8) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_8_0_a3  
        (.A(N_642), .B(N_526), .Y(N_621));
    CFG4 #( .INIT(16'hA0EC) )  
        \clkalign_curr_state_ns_5_0_.un1_RX_CLK_ALIGN_LOAD5_0_1  (.A(
        N_643), .B(N_594_1), .C(N_525), .D(rx_err_Z), .Y(
        un1_RX_CLK_ALIGN_LOAD5_0_1));
    SLE \tapcnt_final[3]  (.D(tapcnt_final_11[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[3]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[23])
        , .D(late_flags_lsb_Z[87]), .FCI(late_found_lsb_126_2_1_co1_17)
        , .S(late_found_lsb_126_2_1_wmux_37_S), .Y(
        late_found_lsb_126_2_1_y0_16), .FCO(
        late_found_lsb_126_2_1_co0_18));
    SLE \late_flags_msb[59]  (.D(late_flags_msb_Z[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[59]));
    CFG4 #( .INIT(16'h04AE) )  \clkalign_curr_state_ns_5_0_.m74_1_1  (
        .A(clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[4]), .C(
        N_19_i), .D(N_30), .Y(m74_1_0));
    SLE \late_flags_lsb[96]  (.D(late_flags_lsb_Z[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[96]));
    SLE \late_flags_lsb[62]  (.D(late_flags_lsb_Z[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[62]));
    SLE \late_flags_msb[75]  (.D(late_flags_msb_Z[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[75]));
    SLE \late_flags_lsb[28]  (.D(late_flags_lsb_Z[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[28]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[22]), .D(early_flags_msb_Z[86]), .FCI(
        early_found_msb_63_2_1_co1_17), .S(
        early_found_msb_63_2_1_wmux_37_S), .Y(
        early_found_msb_63_2_1_y0_16), .FCO(
        early_found_msb_63_2_1_co0_18));
    SLE \early_flags_msb[45]  (.D(early_flags_msb_Z[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[45]));
    SLE \late_flags_lsb[93]  (.D(late_flags_lsb_Z[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[93]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_2 (.A(
        early_found_lsb_63_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[48]), .D(early_flags_lsb_Z[112]), .FCI(
        early_found_lsb_63_2_1_co0_0), .S(
        early_found_lsb_63_2_1_wmux_2_S), .Y(
        early_found_lsb_63_2_1_0_y3), .FCO(
        early_found_lsb_63_2_1_co1_0));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[2]  (.A(
        tapcnt_final_11_iv_1[2]), .B(tapcnt_final_11_iv_0[2]), .Y(
        tapcnt_final_11[2]));
    SLE \sig_tapcnt_final_1[7]  (.D(un3_sig_tapcnt_final_1_cry_7_Z), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[7]));
    SLE \early_flags_lsb[14]  (.D(early_flags_lsb_Z[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[14]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_34 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_63_2_1_co0_16), .S(
        late_found_msb_63_2_1_wmux_34_S), .Y(
        late_found_msb_63_2_1_wmux_34_Y), .FCO(
        late_found_msb_63_2_1_co1_16));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_32 (.A(
        late_found_lsb_126_2_1_y0_14), .B(late_found_lsb_126_2_1_y3_1), 
        .C(late_found_lsb_126_2_1_y1_1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co0_15), .S(
        late_found_lsb_126_2_1_wmux_32_S), .Y(
        late_found_lsb_126_2_1_0_y33), .FCO(
        late_found_lsb_126_2_1_co1_15));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[22])
        , .D(late_flags_msb_Z[86]), .FCI(late_found_msb_63_2_1_co1_17), 
        .S(late_found_msb_63_2_1_wmux_37_S), .Y(
        late_found_msb_63_2_1_y0_16), .FCO(
        late_found_msb_63_2_1_co0_18));
    SLE late_found_lsb_d (.D(late_found_lsb), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(late_found_lsb_d_Z));
    SLE \early_flags_lsb[79]  (.D(early_flags_lsb_Z[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[79]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_nxt_set14_3_i_o3_0  
        (.A(N_525), .B(N_533), .Y(N_549));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[6]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_7_S), 
        .Y(sig_tapcnt_final_2_3_Z[6]));
    SLE \early_flags_msb[70]  (.D(early_flags_msb_Z[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[70]));
    SLE \late_flags_lsb[70]  (.D(late_flags_lsb_Z[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[70]));
    SLE \late_flags_msb[42]  (.D(late_flags_msb_Z[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[42]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_33 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_63_2_1_co1_15), .S(
        early_found_lsb_63_2_1_wmux_33_S), .Y(
        early_found_lsb_63_2_1_wmux_33_Y), .FCO(
        early_found_lsb_63_2_1_co0_16));
    CFG4 #( .INIT(16'h0448) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_i_a2[0]  (.A(
        clkalign_curr_state_Z[4]), .B(N_627), .C(
        clkalign_curr_state_Z[2]), .D(clkalign_curr_state_Z[1]), .Y(
        N_659));
    SLE \late_flags_lsb[105]  (.D(late_flags_lsb_Z[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[105]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[0]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[0]), .D(GND), .FCI(
        emflag_cnt_cry_cy), .S(emflag_cnt_s[0]), .Y(
        emflag_cnt_cry_Y[0]), .FCO(emflag_cnt_cry_Z[0]));
    SLE \early_flags_lsb[54]  (.D(early_flags_lsb_Z[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[54]));
    SLE \late_flags_lsb[88]  (.D(late_flags_lsb_Z[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[88]));
    SLE \tapcnt_final[4]  (.D(tapcnt_final_11[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[4]));
    SLE \early_flags_lsb[11]  (.D(early_flags_lsb_Z[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[11]));
    CFG2 #( .INIT(4'hE) )  early_or_late_found_lsb (.A(
        early_found_lsb_d_Z), .B(late_found_lsb_d_Z), .Y(
        early_or_late_found_lsb_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[19])
        , .D(late_flags_lsb_Z[83]), .FCI(late_found_lsb_126_2_1_co1_11)
        , .S(late_found_lsb_126_2_1_wmux_25_S), .Y(
        late_found_lsb_126_2_1_y0_11), .FCO(
        late_found_lsb_126_2_1_co0_12));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[6]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[6]), .D(GND), .FCI(
        emflag_cnt_cry_Z[5]), .S(emflag_cnt_s[6]), .Y(
        emflag_cnt_cry_Y[6]), .FCO(emflag_cnt_cry_Z[6]));
    SLE \late_flags_msb[32]  (.D(late_flags_msb_Z[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[32]));
    CFG3 #( .INIT(8'h02) )  
        \clkalign_curr_state_ns_5_0_.clk_align_start6_0_a2  (.A(
        clkalign_curr_state_Z[5]), .B(clkalign_curr_state_Z[3]), .C(
        clkalign_curr_state_Z[0]), .Y(N_651));
    SLE \early_flags_lsb[51]  (.D(early_flags_lsb_Z[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[51]));
    SLE \early_flags_lsb[16]  (.D(early_flags_lsb_Z[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[16]));
    SLE \early_flags_msb[108]  (.D(early_flags_msb_Z[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[108]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[16]), .D(early_flags_lsb_Z[80]), .FCI(
        early_found_lsb_63_2_1_0_co1), .S(
        early_found_lsb_63_2_1_wmux_1_S), .Y(
        early_found_lsb_63_2_1_y0_0), .FCO(
        early_found_lsb_63_2_1_co0_0));
    SLE \early_flags_msb[114]  (.D(early_flags_msb_Z[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[114]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[0])
        , .D(early_flags_msb_Z[64]), .FCI(VCC), .S(
        early_found_msb_63_2_1_0_wmux_S), .Y(
        early_found_msb_63_2_1_0_y0), .FCO(
        early_found_msb_63_2_1_0_co0));
    CFG3 #( .INIT(8'hF8) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_14_0  (.A(
        N_653), .B(N_593), .C(clkalign_curr_state_s9_0_a3), .Y(
        un1_clkalign_curr_state_14_0));
    SLE \late_flags_msb[68]  (.D(late_flags_msb_Z[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[68]));
    CFG3 #( .INIT(8'h47) )  \clkalign_curr_state_ns_5_0_.m96_1_1  (.A(
        N_30), .B(clkalign_curr_state_Z[1]), .C(N_78), .Y(m96_1_0));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_26 (.A(
        early_found_lsb_126_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[51]), .D(early_flags_lsb_Z[115]), .FCI(
        early_found_lsb_126_2_1_co0_12), .S(
        early_found_lsb_126_2_1_wmux_26_S), .Y(
        early_found_lsb_126_2_1_y3_1), .FCO(
        early_found_lsb_126_2_1_co1_12));
    SLE \early_flags_msb[95]  (.D(early_flags_msb_Z[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[95]));
    SLE \tapcnt_offset[7]  (.D(tapcnt_offset_s[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[7]));
    CFG4 #( .INIT(16'h74FC) )  \clkalign_curr_state_ns_5_0_.m100  (.A(
        calc_done_Z), .B(clkalign_curr_state_Z[0]), .C(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), .D(N_125_mux), .Y(
        N_101));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_8 (.A(
        late_found_msb_63_2_1_y0_3), .B(late_found_msb_63_2_1_0_y3), 
        .C(late_found_msb_63_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co0_3), .S(
        late_found_msb_63_2_1_wmux_8_S), .Y(late_found_msb_63_2_1_0_y9)
        , .FCO(late_found_msb_63_2_1_co1_3));
    SLE \late_flags_msb[82]  (.D(late_flags_msb_Z[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[82]));
    SLE \early_flags_lsb[56]  (.D(early_flags_lsb_Z[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[56]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[27]), .D(early_flags_lsb_Z[91]), .FCI(
        early_found_lsb_126_2_1_co1_13), .S(
        early_found_lsb_126_2_1_wmux_29_S), .Y(
        early_found_lsb_126_2_1_y0_13), .FCO(
        early_found_lsb_126_2_1_co0_14));
    SLE \late_flags_msb[123]  (.D(late_flags_msb_Z[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[123]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[30]), .D(early_flags_msb_Z[94]), .FCI(
        early_found_msb_63_2_1_co1_19), .S(
        early_found_msb_63_2_1_wmux_41_S), .Y(
        early_found_msb_63_2_1_y0_18), .FCO(
        early_found_msb_63_2_1_co0_20));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_34 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_126_2_1_co0_16), .S(
        early_found_msb_126_2_1_wmux_34_S), .Y(
        early_found_msb_126_2_1_wmux_34_Y), .FCO(
        early_found_msb_126_2_1_co1_16));
    SLE \early_flags_lsb[82]  (.D(early_flags_lsb_Z[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[82]));
    SLE \rst_cnt[3]  (.D(rst_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[3]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_40 (.A(
        early_found_lsb_63_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[46]), .D(early_flags_lsb_Z[110]), .FCI(
        early_found_lsb_63_2_1_co0_19), .S(
        early_found_lsb_63_2_1_wmux_40_S), .Y(
        early_found_lsb_63_2_1_y5_2), .FCO(
        early_found_lsb_63_2_1_co1_19));
    SLE \tapcnt_offset[2]  (.D(tapcnt_offset_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[2]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[6]), 
        .D(late_flags_msb_Z[70]), .FCI(late_found_msb_63_2_1_co1_16), 
        .S(late_found_msb_63_2_1_wmux_35_S), .Y(
        late_found_msb_63_2_1_y0_15), .FCO(
        late_found_msb_63_2_1_co0_17));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_6 
        (.A(early_late_nxt_val_Z[6]), .B(early_late_init_val_Z[6]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_5_Z), 
        .S(early_late_init_nxt_val_status5_cry_6_S), .Y(
        early_late_init_nxt_val_status5_cry_6_Y), .FCO(
        early_late_init_nxt_val_status5_cry_6_Z));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_3 
        (.A(early_late_nxt_val_Z[3]), .B(early_late_init_val_Z[3]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_2_Z), 
        .S(early_late_init_nxt_val_status5_cry_3_S), .Y(
        early_late_init_nxt_val_status5_cry_3_Y), .FCO(
        early_late_init_nxt_val_status5_cry_3_Z));
    CFG3 #( .INIT(8'h27) )  early_found_msb_127_i (.A(emflag_cnt_Z[0]), 
        .B(N_2221), .C(N_2158), .Y(early_found_msb_i));
    CFG2 #( .INIT(4'h8) )  no_early_and_late_found_lsb (.A(
        early_not_found_lsb_d_Z), .B(late_not_found_lsb_d_Z), .Y(
        no_early_and_late_found_lsb_Z));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[3]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[3]), .D(GND), .FCI(
        tap_cnt_cry_Z[2]), .S(tap_cnt_s[3]), .Y(tap_cnt_cry_Y[3]), 
        .FCO(tap_cnt_cry_Z[3]));
    SLE \early_flags_lsb[18]  (.D(early_flags_lsb_Z[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[18]));
    CFG2 #( .INIT(4'h6) )  \clkalign_curr_state_ns_5_0_.m4  (.A(
        clkalign_curr_state_Z[0]), .B(N_125_mux), .Y(N_5));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_12 (.A(
        early_found_msb_126_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[37]), .D(early_flags_msb_Z[101]), .FCI(
        early_found_msb_126_2_1_co0_5), .S(
        early_found_msb_126_2_1_wmux_12_S), .Y(
        early_found_msb_126_2_1_y1_0), .FCO(
        early_found_msb_126_2_1_co1_5));
    SLE \early_flags_msb[17]  (.D(early_flags_msb_Z[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[17]));
    SLE \early_flags_lsb[99]  (.D(early_flags_lsb_Z[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[99]));
    CFG2 #( .INIT(4'h8) )  emflag_cnt_done_0 (.A(emflag_cnt_Z[0]), .B(
        emflag_cnt_Z[7]), .Y(emflag_cnt_done_0_Z));
    SLE \late_flags_msb[127]  (.D(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[127]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_6 (.A(
        late_found_msb_126_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[57]), .D(late_flags_msb_Z[121]), .FCI(
        late_found_msb_126_2_1_co0_2), .S(
        late_found_msb_126_2_1_wmux_6_S), .Y(
        late_found_msb_126_2_1_0_y7), .FCO(
        late_found_msb_126_2_1_co1_2));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[7]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[7]), .D(early_late_start_val_Z[7]), 
        .Y(tapcnt_final_11_iv_0[7]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[26])
        , .D(late_flags_lsb_Z[90]), .FCI(late_found_lsb_63_2_1_co1_13), 
        .S(late_found_lsb_63_2_1_wmux_29_S), .Y(
        late_found_lsb_63_2_1_y0_13), .FCO(
        late_found_lsb_63_2_1_co0_14));
    CFG4 #( .INIT(16'h00F2) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_i_0_RNIUV6P1[0]  (.A(
        N_511_i_1), .B(N_537), .C(wait_cnt_Z[0]), .D(wait_cnt_3_i_0[0])
        , .Y(N_511_i));
    SLE \tapcnt_final[2]  (.D(tapcnt_final_11[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[2]));
    SLE \early_flags_lsb[58]  (.D(early_flags_lsb_Z[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[58]));
    SLE \late_flags_lsb[29]  (.D(late_flags_lsb_Z[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[29]));
    SLE \early_flags_msb[89]  (.D(early_flags_msb_Z[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[89]));
    SLE \late_flags_lsb[7]  (.D(late_flags_lsb_Z[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[7]));
    SLE \early_flags_lsb[39]  (.D(early_flags_lsb_Z[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[39]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_4 (.A(
        early_found_lsb_126_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[41]), .D(early_flags_lsb_Z[105]), .FCI(
        early_found_lsb_126_2_1_co0_1), .S(
        early_found_lsb_126_2_1_wmux_4_S), .Y(
        early_found_lsb_126_2_1_0_y5), .FCO(
        early_found_lsb_126_2_1_co1_1));
    SLE \late_flags_lsb[89]  (.D(late_flags_lsb_Z[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[89]));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[3]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_4_S), 
        .Y(sig_tapcnt_final_1_3_Z[3]));
    SLE \late_flags_lsb[121]  (.D(late_flags_lsb_Z[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[121]));
    SLE \tapcnt_final[0]  (.D(tapcnt_final_11[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[0]));
    SLE \late_flags_msb[92]  (.D(late_flags_msb_Z[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[92]));
    SLE \early_flags_msb[29]  (.D(early_flags_msb_Z[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[29]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[31]), .D(early_flags_msb_Z[95]), .FCI(
        early_found_msb_126_2_1_co1_19), .S(
        early_found_msb_126_2_1_wmux_41_S), .Y(
        early_found_msb_126_2_1_y0_18), .FCO(
        early_found_msb_126_2_1_co0_20));
    CFG3 #( .INIT(8'h01) )  \clkalign_curr_state_ns_5_0_.m9  (.A(
        wait_cnt_Z[2]), .B(wait_cnt_Z[1]), .C(wait_cnt_Z[0]), .Y(
        N_127_mux));
    SLE \late_flags_lsb[67]  (.D(late_flags_lsb_Z[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[67]));
    SLE \early_flags_msb[113]  (.D(early_flags_msb_Z[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[113]));
    SLE \late_flags_lsb[5]  (.D(late_flags_lsb_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[5]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_3 
        (.A(early_late_end_val_Z[3]), .B(early_late_start_val_Z[3]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_2_Z), .S(
        early_late_start_end_val_status5_cry_3_S), .Y(
        early_late_start_end_val_status5_cry_3_Y), .FCO(
        early_late_start_end_val_status5_cry_3_Z));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_30 (.A(
        late_found_msb_126_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[59]), .D(late_flags_msb_Z[123]), .FCI(
        late_found_msb_126_2_1_co0_14), .S(
        late_found_msb_126_2_1_wmux_30_S), .Y(
        late_found_msb_126_2_1_y7_1), .FCO(
        late_found_msb_126_2_1_co1_14));
    SLE \rst_cnt[6]  (.D(rst_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[6]));
    CFG2 #( .INIT(4'h8) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_0_sqmuxa_4_0_a2_0  
        (.A(clkalign_curr_state_RNIJB1J_Y[0]), .B(
        clkalign_curr_state_Z[5]), .Y(N_656));
    SLE \late_flags_msb[28]  (.D(late_flags_msb_Z[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[28]));
    SLE \late_flags_msb[113]  (.D(late_flags_msb_Z[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[113]));
    SLE \emflag_cnt[4]  (.D(emflag_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[4]));
    CFG4 #( .INIT(16'h7351) )  \clkalign_curr_state_ns_5_0_.m62  (.A(
        clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[1]), .C(
        N_61), .D(N_130_mux), .Y(N_63));
    SLE \late_flags_msb[47]  (.D(late_flags_msb_Z[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[47]));
    SLE \early_flags_lsb[47]  (.D(early_flags_lsb_Z[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[47]));
    CFG4 #( .INIT(16'hFFCE) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_1_sqmuxa_5_0  
        (.A(N_643), .B(N_621), .C(N_525), .D(
        un1_clkalign_curr_state_1_sqmuxa_5_0_0), .Y(
        un1_clkalign_curr_state_1_sqmuxa_5_0));
    CFG4 #( .INIT(16'h4073) )  \clkalign_curr_state_ns_5_0_.m57_1_2  (
        .A(clkalign_curr_state_Z[0]), .B(clkalign_curr_state_Z[1]), .C(
        N_55), .D(N_130_mux), .Y(m57_1_2));
    SLE \sig_tapcnt_final_2[2]  (.D(sig_tapcnt_final_2_3_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[2]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_6 (.A(
        early_found_lsb_126_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[57]), .D(early_flags_lsb_Z[121]), .FCI(
        early_found_lsb_126_2_1_co0_2), .S(
        early_found_lsb_126_2_1_wmux_6_S), .Y(
        early_found_lsb_126_2_1_0_y7), .FCO(
        early_found_lsb_126_2_1_co1_2));
    SLE \late_flags_msb[69]  (.D(late_flags_msb_Z[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[69]));
    SLE \sig_tapcnt_final_1[0]  (.D(sig_tapcnt_final_1_3_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[13])
        , .D(late_flags_lsb_Z[77]), .FCI(late_found_lsb_126_2_1_co1_6), 
        .S(late_found_lsb_126_2_1_wmux_15_S), .Y(
        late_found_lsb_126_2_1_y0_7), .FCO(
        late_found_lsb_126_2_1_co0_7));
    SLE \late_flags_lsb[12]  (.D(late_flags_lsb_Z[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[12]));
    SLE \early_flags_msb[14]  (.D(early_flags_msb_Z[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[14]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[5]  (.A(
        tapcnt_final_11_iv_1[5]), .B(tapcnt_final_11_iv_0[5]), .Y(
        tapcnt_final_11[5]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_16 (.A(
        late_found_msb_63_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[44]), .D(late_flags_msb_Z[108]), .FCI(
        late_found_msb_63_2_1_co0_7), .S(
        late_found_msb_63_2_1_wmux_16_S), .Y(
        late_found_msb_63_2_1_y5_0), .FCO(late_found_msb_63_2_1_co1_7));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_3 (.A(
        early_late_end_val_Z[3]), .B(early_late_start_val_Z[3]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_2_Z), .S(
        un3_sig_tapcnt_final_1_cry_3_S), .Y(
        un3_sig_tapcnt_final_1_cry_3_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_3_Z));
    SLE \sig_tapcnt_final_1[1]  (.D(sig_tapcnt_final_1_3_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[1]));
    SLE \late_flags_msb[117]  (.D(late_flags_msb_Z[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[117]));
    SLE \early_late_start_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[1]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_28 (.A(
        early_found_lsb_126_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[43]), .D(early_flags_lsb_Z[107]), .FCI(
        early_found_lsb_126_2_1_co0_13), .S(
        early_found_lsb_126_2_1_wmux_28_S), .Y(
        early_found_lsb_126_2_1_y5_1), .FCO(
        early_found_lsb_126_2_1_co1_13));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_30 (.A(
        early_found_lsb_126_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[59]), .D(early_flags_lsb_Z[123]), .FCI(
        early_found_lsb_126_2_1_co0_14), .S(
        early_found_lsb_126_2_1_wmux_30_S), .Y(
        early_found_lsb_126_2_1_y7_1), .FCO(
        early_found_lsb_126_2_1_co1_14));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_30 (.A(
        late_found_msb_63_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[58]), .D(late_flags_msb_Z[122]), .FCI(
        late_found_msb_63_2_1_co0_14), .S(
        late_found_msb_63_2_1_wmux_30_S), .Y(
        late_found_msb_63_2_1_y7_1), .FCO(late_found_msb_63_2_1_co1_14)
        );
    SLE \early_flags_lsb[85]  (.D(early_flags_lsb_Z[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[85]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_36 (.A(
        late_found_lsb_63_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[38]), .D(late_flags_lsb_Z[102]), .FCI(
        late_found_lsb_63_2_1_co0_17), .S(
        late_found_lsb_63_2_1_wmux_36_S), .Y(
        late_found_lsb_63_2_1_y1_2), .FCO(late_found_lsb_63_2_1_co1_17)
        );
    CFG4 #( .INIT(16'h31B9) )  \clkalign_curr_state_ns_5_0_.m114_2_1  
        (.A(clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), 
        .C(N_137_mux), .D(clkalign_curr_state_Z[4]), .Y(m114_2_1));
    SLE \early_flags_lsb[63]  (.D(early_flags_lsb_Z[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[63]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[2]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[2]), .D(GND), .FCI(
        emflag_cnt_cry_Z[1]), .S(emflag_cnt_s[2]), .Y(
        emflag_cnt_cry_Y[2]), .FCO(emflag_cnt_cry_Z[2]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[19])
        , .D(late_flags_msb_Z[83]), .FCI(late_found_msb_126_2_1_co1_11)
        , .S(late_found_msb_126_2_1_wmux_25_S), .Y(
        late_found_msb_126_2_1_y0_11), .FCO(
        late_found_msb_126_2_1_co0_12));
    SLE \late_flags_msb[37]  (.D(late_flags_msb_Z[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[37]));
    CFG3 #( .INIT(8'hED) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3[1]  (.A(N_546), .B(
        N_540), .C(wait_cnt_Z[1]), .Y(wait_cnt_3[1]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_12 (.A(
        early_found_lsb_126_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[37]), .D(early_flags_lsb_Z[101]), .FCI(
        early_found_lsb_126_2_1_co0_5), .S(
        early_found_lsb_126_2_1_wmux_12_S), .Y(
        early_found_lsb_126_2_1_y1_0), .FCO(
        early_found_lsb_126_2_1_co1_5));
    CFG3 #( .INIT(8'h02) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s9_0_a3  (.A(
        N_2979), .B(N_525), .C(N_533), .Y(clkalign_curr_state_s9_0_a3));
    CFG4 #( .INIT(16'hFFFE) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_o2[1]  (.A(N_537), .B(
        wait_cnt_Z[0]), .C(clkalign_curr_state_Z[3]), .D(
        clkalign_curr_state_Z[0]), .Y(N_546));
    SLE \late_flags_lsb[64]  (.D(late_flags_lsb_Z[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[64]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[6]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[6]), .D(early_late_start_val_Z[6]), 
        .Y(tapcnt_final_11_iv_0[6]));
    SLE \early_flags_msb[11]  (.D(early_flags_msb_Z[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[11]));
    SLE \early_flags_lsb[126]  (.D(early_flags_lsb_Z[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[126]));
    CFG4 #( .INIT(16'h5D00) )  \clkalign_curr_state_ns_5_0_.m108  (.A(
        clkalign_curr_state_Z[4]), .B(early_or_late_found_Z), .C(
        emflag_cnt_done_d_Z), .D(clkalign_curr_state_Z[0]), .Y(N_109));
    CFG4 #( .INIT(16'h0001) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_end_set12_3_i_a3  
        (.A(emflag_cnt_done_d_Z), .B(clkalign_curr_state_Z[3]), .C(
        early_or_late_found_Z), .D(no_early_and_late_found_Z), .Y(
        N_619));
    CFG2 #( .INIT(4'h1) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s5_0_a2  (.A(
        clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[5]), .Y(
        N_627));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[2])
        , .D(early_flags_msb_Z[66]), .FCI(
        early_found_msb_63_2_1_co1_10), .S(
        early_found_msb_63_2_1_wmux_23_S), .Y(
        early_found_msb_63_2_1_y0_10), .FCO(
        early_found_msb_63_2_1_co0_11));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_12 (.A(
        late_found_lsb_63_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[36]), .D(late_flags_lsb_Z[100]), .FCI(
        late_found_lsb_63_2_1_co0_5), .S(
        late_found_lsb_63_2_1_wmux_12_S), .Y(
        late_found_lsb_63_2_1_y1_0), .FCO(late_found_lsb_63_2_1_co1_5));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_6 
        (.A(early_late_end_val_Z[6]), .B(early_late_start_val_Z[6]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_5_Z), .S(
        early_late_start_end_val_status5_cry_6_S), .Y(
        early_late_start_end_val_status5_cry_6_Y), .FCO(
        early_late_start_end_val_status5_cry_6_Z));
    SLE \late_flags_msb[87]  (.D(late_flags_msb_Z[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[87]));
    SLE \late_flags_msb[44]  (.D(late_flags_msb_Z[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[44]));
    SLE \tap_cnt[5]  (.D(tap_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[5]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_26 (.A(
        late_found_msb_63_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[50]), .D(late_flags_msb_Z[114]), .FCI(
        late_found_msb_63_2_1_co0_12), .S(
        late_found_msb_63_2_1_wmux_26_S), .Y(
        late_found_msb_63_2_1_y3_1), .FCO(late_found_msb_63_2_1_co1_12)
        );
    SLE \early_flags_msb[16]  (.D(early_flags_msb_Z[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[16]));
    SLE \late_flags_lsb[111]  (.D(late_flags_lsb_Z[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[111]));
    SLE \early_flags_lsb[23]  (.D(early_flags_lsb_Z[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[23]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_42 (.A(
        late_found_msb_126_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[63]), .D(late_flags_msb_Z[127]), .FCI(
        late_found_msb_126_2_1_co0_20), .S(
        late_found_msb_126_2_1_wmux_42_S), .Y(
        late_found_msb_126_2_1_y7_2), .FCO(
        late_found_msb_126_2_1_co1_20));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[20]), .D(early_flags_msb_Z[84]), .FCI(
        early_found_msb_63_2_1_co1_5), .S(
        early_found_msb_63_2_1_wmux_13_S), .Y(
        early_found_msb_63_2_1_y0_6), .FCO(
        early_found_msb_63_2_1_co0_6));
    CFG3 #( .INIT(8'hEA) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_1_0  (.A(
        clkalign_curr_state_s9_0_a3), .B(
        un1_clkalign_curr_state_1_0_a3_0), .C(N_627), .Y(
        un1_clkalign_curr_state_1_0));
    SLE tapcnt_final_2_status (.D(sig_tapcnt_final_210_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_final_2_status_Z));
    CFG4 #( .INIT(16'h0001) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state63_NE_i  (.A(
        clkalign_curr_state63_NE_0), .B(clkalign_curr_state63_NE_3), 
        .C(clkalign_curr_state63_NE_2), .D(clkalign_curr_state63_NE_1), 
        .Y(clkalign_curr_state63));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_8 (.A(
        early_found_lsb_126_2_1_y0_3), .B(early_found_lsb_126_2_1_0_y3)
        , .C(early_found_lsb_126_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_126_2_1_co0_3), .S(
        early_found_lsb_126_2_1_wmux_8_S), .Y(
        early_found_lsb_126_2_1_0_y9), .FCO(
        early_found_lsb_126_2_1_co1_3));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_2 (.A(
        early_found_lsb_126_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[49]), .D(early_flags_lsb_Z[113]), .FCI(
        early_found_lsb_126_2_1_co0_0), .S(
        early_found_lsb_126_2_1_wmux_2_S), .Y(
        early_found_lsb_126_2_1_0_y3), .FCO(
        early_found_lsb_126_2_1_co1_0));
    SLE \tapcnt_final[7]  (.D(tapcnt_final_11[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[7]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_42 (.A(
        late_found_msb_63_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[62]), .D(late_flags_msb_Z[126]), .FCI(
        late_found_msb_63_2_1_co0_20), .S(
        late_found_msb_63_2_1_wmux_42_S), .Y(
        late_found_msb_63_2_1_y7_2), .FCO(late_found_msb_63_2_1_co1_20)
        );
    SLE \late_flags_lsb[90]  (.D(late_flags_lsb_Z[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[90]));
    SLE \early_flags_lsb[70]  (.D(early_flags_lsb_Z[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[70]));
    CFG3 #( .INIT(8'hB8) )  \clkalign_curr_state_ns_5_0_.m115  (.A(
        N_115), .B(clkalign_curr_state_Z[3]), .C(N_132_mux), .Y(N_116));
    SLE early_late_end_set (.D(clkalign_curr_state_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(N_515_i), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_late_end_set_Z));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_21 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_126_2_1_co1_9), .S(
        early_found_msb_126_2_1_wmux_21_S), .Y(
        early_found_msb_126_2_1_wmux_21_Y), .FCO(
        early_found_msb_126_2_1_co0_10));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[4]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[4]), .D(GND), .FCI(
        emflag_cnt_cry_Z[3]), .S(emflag_cnt_s[4]), .Y(
        emflag_cnt_cry_Y[4]), .FCO(emflag_cnt_cry_Z[4]));
    SLE \early_flags_lsb[106]  (.D(early_flags_lsb_Z[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[106]));
    SLE \early_flags_lsb[44]  (.D(early_flags_lsb_Z[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[44]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[5]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[5]), .D(GND), .FCI(
        emflag_cnt_cry_Z[4]), .S(emflag_cnt_s[5]), .Y(
        emflag_cnt_cry_Y[5]), .FCO(emflag_cnt_cry_Z[5]));
    SLE \late_flags_msb[34]  (.D(late_flags_msb_Z[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[34]));
    CFG4 #( .INIT(16'h5C50) )  \clkalign_curr_state_ns_5_0_.m11  (.A(
        N_125_mux), .B(PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), .C(
        clkalign_curr_state_Z[0]), .D(N_127_mux), .Y(N_12));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_cry[1]  (.A(VCC), .B(
        timeout_cnt_Z[1]), .C(GND), .D(GND), .FCI(
        timeout_cnt_s_1134_FCO), .S(timeout_cnt_s[1]), .Y(
        timeout_cnt_cry_Y[1]), .FCO(timeout_cnt_cry_Z[1]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[2]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[2]), .D(early_late_init_val_Z[2]), .Y(
        tapcnt_final_11_iv_1[2]));
    SLE \early_flags_msb[18]  (.D(early_flags_msb_Z[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[18]));
    SLE \late_flags_msb[100]  (.D(late_flags_msb_Z[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[100]));
    SLE \rst_cnt[1]  (.D(rst_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[1]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_22 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_126_2_1_co0_10), .S(
        late_found_msb_126_2_1_wmux_22_S), .Y(
        late_found_msb_126_2_1_wmux_22_Y), .FCO(
        late_found_msb_126_2_1_co1_10));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[9]), 
        .D(late_flags_lsb_Z[73]), .FCI(late_found_lsb_126_2_1_co1_0), 
        .S(late_found_lsb_126_2_1_wmux_3_S), .Y(
        late_found_lsb_126_2_1_y0_1), .FCO(
        late_found_lsb_126_2_1_co0_1));
    SLE \late_flags_msb[29]  (.D(late_flags_msb_Z[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[29]));
    CFG4 #( .INIT(16'h0001) )  \clkalign_curr_state_ns_5_0_.m77  (.A(
        wait_cnt_Z[0]), .B(clkalign_curr_state_Z[0]), .C(wait_cnt_Z[2])
        , .D(wait_cnt_Z[1]), .Y(N_78));
    SLE \late_flags_msb[84]  (.D(late_flags_msb_Z[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[84]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_40 (.A(
        early_found_msb_63_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[46]), .D(early_flags_msb_Z[110]), .FCI(
        early_found_msb_63_2_1_co0_19), .S(
        early_found_msb_63_2_1_wmux_40_S), .Y(
        early_found_msb_63_2_1_y5_2), .FCO(
        early_found_msb_63_2_1_co1_19));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_28 (.A(
        late_found_msb_126_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[43]), .D(late_flags_msb_Z[107]), .FCI(
        late_found_msb_126_2_1_co0_13), .S(
        late_found_msb_126_2_1_wmux_28_S), .Y(
        late_found_msb_126_2_1_y5_1), .FCO(
        late_found_msb_126_2_1_co1_13));
    SLE \early_flags_lsb[12]  (.D(early_flags_lsb_Z[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[12]));
    SLE \early_flags_lsb[41]  (.D(early_flags_lsb_Z[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[41]));
    SLE \early_late_init_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[4]));
    SLE late_found_msb_d (.D(late_found_msb), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(late_found_msb_d_Z));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_126_2_1_wmux_7 (.A(
        late_found_msb_126_2_1_0_y7), .B(late_found_msb_126_2_1_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co1_2), .S(
        late_found_msb_126_2_1_wmux_7_S), .Y(
        late_found_msb_126_2_1_y0_3), .FCO(
        late_found_msb_126_2_1_co0_3));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_14 (.A(
        late_found_lsb_63_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[52]), .D(late_flags_lsb_Z[116]), .FCI(
        late_found_lsb_63_2_1_co0_6), .S(
        late_found_lsb_63_2_1_wmux_14_S), .Y(
        late_found_lsb_63_2_1_y3_0), .FCO(late_found_lsb_63_2_1_co1_6));
    SLE \early_flags_msb[0]  (.D(early_flags_msb_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[0]));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_1 (.A(
        early_late_end_val_Z[1]), .B(early_late_start_val_Z[1]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_0_Z), .S(
        un3_sig_tapcnt_final_1_cry_1_S), .Y(
        un3_sig_tapcnt_final_1_cry_1_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_1_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[28])
        , .D(late_flags_lsb_Z[92]), .FCI(late_found_lsb_63_2_1_co1_7), 
        .S(late_found_lsb_63_2_1_wmux_17_S), .Y(
        late_found_lsb_63_2_1_y0_8), .FCO(late_found_lsb_63_2_1_co0_8));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[21]), .D(early_flags_msb_Z[85]), .FCI(
        early_found_msb_126_2_1_co1_5), .S(
        early_found_msb_126_2_1_wmux_13_S), .Y(
        early_found_msb_126_2_1_y0_6), .FCO(
        early_found_msb_126_2_1_co0_6));
    SLE \late_flags_msb[101]  (.D(late_flags_msb_Z[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[101]));
    ARI1 #( .INIT(20'h44400) )  \emflag_cnt_cry_cy[0]  (.A(VCC), .B(
        N_2979), .C(clkalign_curr_state_Z[0]), .D(GND), .FCI(VCC), .S(
        emflag_cnt_cry_cy_S[0]), .Y(emflag_cnt_cry_cy_Y[0]), .FCO(
        emflag_cnt_cry_cy));
    SLE \late_flags_msb[97]  (.D(late_flags_msb_Z[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[97]));
    SLE \early_flags_msb[5]  (.D(early_flags_msb_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[5]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_28 (.A(
        late_found_lsb_126_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[43]), .D(late_flags_lsb_Z[107]), .FCI(
        late_found_lsb_126_2_1_co0_13), .S(
        late_found_lsb_126_2_1_wmux_28_S), .Y(
        late_found_lsb_126_2_1_y5_1), .FCO(
        late_found_lsb_126_2_1_co1_13));
    SLE \early_flags_lsb[8]  (.D(early_flags_lsb_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[8]));
    SLE early_late_start_end_val_status (.D(
        early_late_start_end_val_status5), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_late_start_end_val_status_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_63_2_1_wmux_31 (.A(
        early_found_lsb_63_2_1_y7_1), .B(early_found_lsb_63_2_1_y5_1), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co1_14), .S(
        early_found_lsb_63_2_1_wmux_31_S), .Y(
        early_found_lsb_63_2_1_y0_14), .FCO(
        early_found_lsb_63_2_1_co0_15));
    SLE \early_flags_lsb[52]  (.D(early_flags_lsb_Z[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[52]));
    SLE \late_flags_lsb[56]  (.D(late_flags_lsb_Z[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[56]));
    SLE \late_flags_lsb[127]  (.D(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[127]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_0 
        (.A(early_late_end_val_Z[0]), .B(early_late_start_val_Z[0]), 
        .C(GND), .D(GND), .FCI(GND), .S(
        early_late_start_end_val_status5_cry_0_S), .Y(
        early_late_start_end_val_status5_cry_0_Y), .FCO(
        early_late_start_end_val_status5_cry_0_Z));
    SLE \early_flags_lsb[46]  (.D(early_flags_lsb_Z[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[46]));
    SLE \late_flags_lsb[42]  (.D(late_flags_lsb_Z[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[42]));
    SLE \late_flags_lsb[53]  (.D(late_flags_lsb_Z[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[53]));
    SLE \wait_cnt[0]  (.D(N_511_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(wait_cnt_Z[0]));
    CFG4 #( .INIT(16'h0004) )  \clkalign_curr_state_ns_5_0_.m122_0_0  
        (.A(clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[4]), 
        .C(clkalign_curr_state_Z[3]), .D(clkalign_curr_state_Z[2]), .Y(
        m122_0_0));
    SLE \early_flags_msb[53]  (.D(early_flags_msb_Z[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[53]));
    SLE \clkalign_curr_state[0]  (.D(N_40_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(clkalign_curr_state_Z[0]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_44 (.A(
        late_found_msb_63_2_1_y0_19), .B(late_found_msb_63_2_1_y3_2), 
        .C(late_found_msb_63_2_1_y1_2), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co0_21), .S(
        late_found_msb_63_2_1_wmux_44_S), .Y(
        late_found_msb_63_2_1_0_y45), .FCO(
        late_found_msb_63_2_1_co1_21));
    SLE \late_flags_msb[7]  (.D(late_flags_msb_Z[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[7]));
    SLE \late_flags_lsb[78]  (.D(late_flags_lsb_Z[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[78]));
    SLE \early_late_nxt_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[4]));
    CFG3 #( .INIT(8'hEA) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_1_sqmuxa_5_0_0  
        (.A(clkalign_curr_state_1_sqmuxa_1), .B(
        clkalign_curr_state_RNIJB1J_Y[0]), .C(N_657), .Y(
        un1_clkalign_curr_state_1_sqmuxa_5_0_0));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_63_2_1_wmux_19 (.A(
        late_found_msb_63_2_1_y7_0), .B(late_found_msb_63_2_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co1_8), .S(
        late_found_msb_63_2_1_wmux_19_S), .Y(
        late_found_msb_63_2_1_y0_9), .FCO(late_found_msb_63_2_1_co0_9));
    SLE \tapcnt_offset[3]  (.D(tapcnt_offset_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[3]));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_6 (.A(
        early_late_end_val_Z[6]), .B(early_late_start_val_Z[6]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_5_Z), .S(
        un3_sig_tapcnt_final_1_cry_6_S), .Y(
        un3_sig_tapcnt_final_1_cry_6_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_6_Z));
    SLE \early_flags_msb[77]  (.D(early_flags_msb_Z[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[77]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[1]  (.A(
        tapcnt_final_11_iv_1[1]), .B(tapcnt_final_11_iv_0[1]), .Y(
        tapcnt_final_11[1]));
    SLE \timeout_cnt[6]  (.D(timeout_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[6]));
    SLE \tap_cnt[1]  (.D(tap_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[1]));
    SLE \late_flags_lsb[17]  (.D(late_flags_lsb_Z[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[17]));
    SLE \early_flags_lsb[90]  (.D(early_flags_lsb_Z[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[90]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[14])
        , .D(late_flags_lsb_Z[78]), .FCI(late_found_lsb_63_2_1_co1_18), 
        .S(late_found_lsb_63_2_1_wmux_39_S), .Y(
        late_found_lsb_63_2_1_y0_17), .FCO(
        late_found_lsb_63_2_1_co0_19));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[13])
        , .D(late_flags_msb_Z[77]), .FCI(late_found_msb_126_2_1_co1_6), 
        .S(late_found_msb_126_2_1_wmux_15_S), .Y(
        late_found_msb_126_2_1_y0_7), .FCO(
        late_found_msb_126_2_1_co0_7));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[0])
        , .D(early_flags_lsb_Z[64]), .FCI(VCC), .S(
        early_found_lsb_63_2_1_0_wmux_S), .Y(
        early_found_lsb_63_2_1_0_y0), .FCO(
        early_found_lsb_63_2_1_0_co0));
    CFG3 #( .INIT(8'hC5) )  \clkalign_curr_state_ns_5_0_.m24  (.A(N_17)
        , .B(N_3109_mux), .C(clkalign_curr_state_Z[3]), .Y(N_25));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_63_2_1_wmux_7 (.A(
        late_found_msb_63_2_1_0_y7), .B(late_found_msb_63_2_1_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co1_2), .S(
        late_found_msb_63_2_1_wmux_7_S), .Y(late_found_msb_63_2_1_y0_3)
        , .FCO(late_found_msb_63_2_1_co0_3));
    SLE \early_flags_lsb[115]  (.D(early_flags_lsb_Z[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[115]));
    SLE clk_align_done (.D(clk_align_start6), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_internal_rst_en_2_0), 
        .ALn(current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(clk_align_done_Z));
    SLE \sig_tapcnt_final_1[3]  (.D(sig_tapcnt_final_1_3_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[3]));
    SLE \early_flags_lsb[48]  (.D(early_flags_lsb_Z[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[48]));
    SLE \early_flags_lsb[120]  (.D(early_flags_lsb_Z[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[120]));
    SLE \late_flags_msb[94]  (.D(late_flags_msb_Z[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[94]));
    SLE \late_flags_lsb[32]  (.D(late_flags_lsb_Z[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[32]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_33 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_63_2_1_co1_15), .S(
        early_found_msb_63_2_1_wmux_33_S), .Y(
        early_found_msb_63_2_1_wmux_33_Y), .FCO(
        early_found_msb_63_2_1_co0_16));
    SLE \late_flags_msb[105]  (.D(late_flags_msb_Z[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[105]));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_cry[3]  (.A(VCC), .B(
        timeout_cnt_Z[3]), .C(GND), .D(GND), .FCI(timeout_cnt_cry_Z[2])
        , .S(timeout_cnt_s[3]), .Y(timeout_cnt_cry_Y[3]), .FCO(
        timeout_cnt_cry_Z[3]));
    SLE \early_flags_msb[80]  (.D(early_flags_msb_Z[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[80]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[26])
        , .D(late_flags_msb_Z[90]), .FCI(late_found_msb_63_2_1_co1_13), 
        .S(late_found_msb_63_2_1_wmux_29_S), .Y(
        late_found_msb_63_2_1_y0_13), .FCO(
        late_found_msb_63_2_1_co0_14));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[12])
        , .D(late_flags_lsb_Z[76]), .FCI(late_found_lsb_63_2_1_co1_6), 
        .S(late_found_lsb_63_2_1_wmux_15_S), .Y(
        late_found_lsb_63_2_1_y0_7), .FCO(late_found_lsb_63_2_1_co0_7));
    SLE \early_late_nxt_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[3]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_11_0  (.A(
        N_585_i), .B(N_634_i), .Y(un1_clkalign_curr_state_11_0));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_4 
        (.A(early_late_nxt_val_Z[4]), .B(early_late_init_val_Z[4]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_3_Z), 
        .S(early_late_init_nxt_val_status5_cry_4_S), .Y(
        early_late_init_nxt_val_status5_cry_4_Y), .FCO(
        early_late_init_nxt_val_status5_cry_4_Z));
    CFG3 #( .INIT(8'h08) )  \clkalign_curr_state_ns_5_0_.m60  (.A(
        early_or_late_found_Z), .B(clkalign_curr_state_Z[0]), .C(
        emflag_cnt_done_d_Z), .Y(N_61));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_44 (.A(
        early_found_lsb_63_2_1_y0_19), .B(early_found_lsb_63_2_1_y3_2), 
        .C(early_found_lsb_63_2_1_y1_2), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co0_21), .S(
        early_found_lsb_63_2_1_wmux_44_S), .Y(
        early_found_lsb_63_2_1_0_y45), .FCO(
        early_found_lsb_63_2_1_co1_21));
    SLE \early_flags_lsb[30]  (.D(early_flags_lsb_Z[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[30]));
    CFG2 #( .INIT(4'h8) )  \clkalign_curr_state_ns_5_0_.m31  (.A(
        N_19_i), .B(clkalign_curr_state_Z[4]), .Y(N_32_i));
    SLE \early_flags_msb[122]  (.D(early_flags_msb_Z[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[122]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[24])
        , .D(late_flags_msb_Z[88]), .FCI(late_found_msb_63_2_1_co1_1), 
        .S(late_found_msb_63_2_1_wmux_5_S), .Y(
        late_found_msb_63_2_1_y0_2), .FCO(late_found_msb_63_2_1_co0_2));
    SLE \early_flags_msb[20]  (.D(early_flags_msb_Z[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[20]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[3]  (.A(
        tapcnt_final_11_iv_1[3]), .B(tapcnt_final_11_iv_0[3]), .Y(
        tapcnt_final_11[3]));
    CFG2 #( .INIT(4'h7) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_0_sqmuxa_4_0_o2  
        (.A(clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[1]), 
        .Y(N_523));
    SLE \early_flags_lsb[123]  (.D(early_flags_lsb_Z[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[123]));
    SLE \early_flags_lsb[100]  (.D(early_flags_lsb_Z[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[100]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[31])
        , .D(late_flags_lsb_Z[95]), .FCI(late_found_lsb_126_2_1_co1_19)
        , .S(late_found_lsb_126_2_1_wmux_41_S), .Y(
        late_found_lsb_126_2_1_y0_18), .FCO(
        late_found_lsb_126_2_1_co0_20));
    SLE \late_flags_lsb[14]  (.D(late_flags_lsb_Z[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[14]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[4]  (.A(
        tapcnt_final_11_iv_1[4]), .B(tapcnt_final_11_iv_0[4]), .Y(
        tapcnt_final_11[4]));
    SLE \sig_tapcnt_final_1[6]  (.D(sig_tapcnt_final_1_3_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[6]));
    SLE \late_flags_lsb[117]  (.D(late_flags_lsb_Z[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[117]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_36 (.A(
        early_found_msb_126_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[39]), .D(early_flags_msb_Z[103]), .FCI(
        early_found_msb_126_2_1_co0_17), .S(
        early_found_msb_126_2_1_wmux_36_S), .Y(
        early_found_msb_126_2_1_y1_2), .FCO(
        early_found_msb_126_2_1_co1_17));
    CFG2 #( .INIT(4'h4) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_13_0_0_974_a3  
        (.A(clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[2]), 
        .Y(N_2979));
    SLE \early_flags_msb[39]  (.D(early_flags_msb_Z[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[39]));
    SLE \early_flags_lsb[15]  (.D(early_flags_lsb_Z[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[15]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_38 (.A(
        late_found_msb_63_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[54]), .D(late_flags_msb_Z[118]), .FCI(
        late_found_msb_63_2_1_co0_18), .S(
        late_found_msb_63_2_1_wmux_38_S), .Y(
        late_found_msb_63_2_1_y3_2), .FCO(late_found_msb_63_2_1_co1_18)
        );
    SLE \clkalign_curr_state[2]  (.D(clkalign_curr_state_ns[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(clkalign_curr_state_Z[2]));
    SLE \early_flags_msb[6]  (.D(early_flags_msb_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[6]));
    SLE \early_flags_lsb[3]  (.D(early_flags_lsb_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[3]));
    SLE \early_flags_msb[74]  (.D(early_flags_msb_Z[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[74]));
    SLE \tapcnt_offset[4]  (.D(tapcnt_offset_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[4]));
    SLE \early_late_start_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[4]));
    SLE \timeout_cnt[0]  (.D(timeout_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_12 (.A(
        late_found_msb_126_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[37]), .D(late_flags_msb_Z[101]), .FCI(
        late_found_msb_126_2_1_co0_5), .S(
        late_found_msb_126_2_1_wmux_12_S), .Y(
        late_found_msb_126_2_1_y1_0), .FCO(
        late_found_msb_126_2_1_co1_5));
    SLE \early_flags_msb[102]  (.D(early_flags_msb_Z[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[102]));
    SLE \early_flags_lsb[55]  (.D(early_flags_lsb_Z[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[55]));
    ARI1 #( .INIT(20'h0EA4A) )  late_found_lsb_63_2_1_wmux_9 (.A(
        late_found_lsb_63_2_1_0_y45), .B(late_found_lsb_63_2_1_y0_4), 
        .C(late_found_lsb_63_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        late_found_lsb_63_2_1_co1_3), .S(
        late_found_lsb_63_2_1_wmux_9_S), .Y(N_2031), .FCO(
        late_found_lsb_63_2_1_co0_4));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_18 (.A(
        late_found_msb_126_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[61]), .D(late_flags_msb_Z[125]), .FCI(
        late_found_msb_126_2_1_co0_8), .S(
        late_found_msb_126_2_1_wmux_18_S), .Y(
        late_found_msb_126_2_1_y7_0), .FCO(
        late_found_msb_126_2_1_co1_8));
    SLE \early_flags_lsb[103]  (.D(early_flags_lsb_Z[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[103]));
    SLE \late_flags_lsb[61]  (.D(late_flags_lsb_Z[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[61]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_5 
        (.A(early_late_end_val_Z[5]), .B(early_late_start_val_Z[5]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_4_Z), .S(
        early_late_start_end_val_status5_cry_5_S), .Y(
        early_late_start_end_val_status5_cry_5_Y), .FCO(
        early_late_start_end_val_status5_cry_5_Z));
    SLE \late_flags_lsb[79]  (.D(late_flags_lsb_Z[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[79]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_21 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_126_2_1_co1_9), .S(
        late_found_lsb_126_2_1_wmux_21_S), .Y(
        late_found_lsb_126_2_1_wmux_21_Y), .FCO(
        late_found_lsb_126_2_1_co0_10));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[0]  (.A(
        tapcnt_final_11_iv_1[0]), .B(tapcnt_final_11_iv_0[0]), .Y(
        tapcnt_final_11[0]));
    CFG4 #( .INIT(16'h4F0F) )  \clkalign_curr_state_ns_5_0_.m107  (.A(
        clkalign_curr_state_Z[0]), .B(clkalign_curr_state_Z[2]), .C(
        clkalign_curr_state_Z[4]), .D(clkalign_curr_state_Z[1]), .Y(
        N_132_mux));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_0 (.A(
        early_found_msb_63_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[32]), .D(early_flags_msb_Z[96]), .FCI(
        early_found_msb_63_2_1_0_co0), .S(
        early_found_msb_63_2_1_wmux_0_S), .Y(
        early_found_msb_63_2_1_0_y1), .FCO(
        early_found_msb_63_2_1_0_co1));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_18 (.A(
        late_found_lsb_126_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[61]), .D(late_flags_lsb_Z[125]), .FCI(
        late_found_lsb_126_2_1_co0_8), .S(
        late_found_lsb_126_2_1_wmux_18_S), .Y(
        late_found_lsb_126_2_1_y7_0), .FCO(
        late_found_lsb_126_2_1_co1_8));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_22 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_63_2_1_co0_10), .S(
        late_found_lsb_63_2_1_wmux_22_S), .Y(
        late_found_lsb_63_2_1_wmux_22_Y), .FCO(
        late_found_lsb_63_2_1_co1_10));
    CFG2 #( .INIT(4'h1) )  
        \clkalign_curr_state_ns_5_0_.emflag_cnt10_i_a2  (.A(N_523), .B(
        clkalign_curr_state_Z[2]), .Y(N_657));
    SLE \early_flags_msb[71]  (.D(early_flags_msb_Z[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[71]));
    SLE \late_flags_msb[52]  (.D(late_flags_msb_Z[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[52]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[8]  (.A(VCC), .B(
        rst_cnt_Z[8]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[7]), .S(
        rst_cnt_s[8]), .Y(rst_cnt_cry_Y[8]), .FCO(rst_cnt_cry_Z[8]));
    SLE \late_flags_msb[41]  (.D(late_flags_msb_Z[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[41]));
    SLE \late_flags_lsb[65]  (.D(late_flags_lsb_Z[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[65]));
    SLE \late_flags_lsb[47]  (.D(late_flags_lsb_Z[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[47]));
    SLE RX_CLK_ALIGN_LOAD (.D(N_2935_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_RX_CLK_ALIGN_LOAD5_0)
        , .ALn(current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD));
    SLE \early_flags_msb[12]  (.D(early_flags_msb_Z[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[12]));
    CFG2 #( .INIT(4'hD) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_nxt_set14_3_i_o2  
        (.A(clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[5]), 
        .Y(N_533));
    SLE \early_flags_msb[76]  (.D(early_flags_msb_Z[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[76]));
    SLE \late_flags_msb[16]  (.D(late_flags_msb_Z[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[16]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[11]), .D(early_flags_msb_Z[75]), .FCI(
        early_found_msb_126_2_1_co1_12), .S(
        early_found_msb_126_2_1_wmux_27_S), .Y(
        early_found_msb_126_2_1_y0_12), .FCO(
        early_found_msb_126_2_1_co0_13));
    SLE \late_flags_msb[13]  (.D(late_flags_msb_Z[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[13]));
    SLE \late_flags_msb[45]  (.D(late_flags_msb_Z[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[45]));
    CFG3 #( .INIT(8'hD8) )  early_or_late_found (.A(emflag_cnt_Z[7]), 
        .B(early_or_late_found_msb_d_Z), .C(
        early_or_late_found_lsb_d_Z), .Y(early_or_late_found_Z));
    SLE \early_flags_lsb[1]  (.D(early_flags_lsb_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[1]));
    SLE \early_flags_msb[126]  (.D(early_flags_msb_Z[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[126]));
    SLE \late_flags_msb[104]  (.D(late_flags_msb_Z[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[104]));
    ARI1 #( .INIT(20'h0CEC2) )  late_found_lsb_63_2_1_wmux_10 (.A(
        late_found_lsb_63_2_1_0_y21), .B(late_found_lsb_63_2_1_0_y9), 
        .C(emflag_cnt_Z[2]), .D(emflag_cnt_Z[1]), .FCI(
        late_found_lsb_63_2_1_co0_4), .S(
        late_found_lsb_63_2_1_wmux_10_S), .Y(
        late_found_lsb_63_2_1_y0_4), .FCO(late_found_lsb_63_2_1_co1_4));
    SLE \late_flags_lsb[126]  (.D(late_flags_lsb_Z[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[126]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_22 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_63_2_1_co0_10), .S(
        early_found_lsb_63_2_1_wmux_22_S), .Y(
        early_found_lsb_63_2_1_wmux_22_Y), .FCO(
        early_found_lsb_63_2_1_co1_10));
    SLE \late_flags_msb[31]  (.D(late_flags_msb_Z[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[31]));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[4]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[4]), .D(GND), .FCI(
        tap_cnt_cry_Z[3]), .S(tap_cnt_s[4]), .Y(tap_cnt_cry_Y[4]), 
        .FCO(tap_cnt_cry_Z[4]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[2]  (.A(VCC), .B(
        rst_cnt_Z[2]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[1]), .S(
        rst_cnt_s[2]), .Y(rst_cnt_cry_Y[2]), .FCO(rst_cnt_cry_Z[2]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_2 
        (.A(early_late_end_val_Z[2]), .B(early_late_start_val_Z[2]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_1_Z), .S(
        early_late_start_end_val_status5_cry_2_S), .Y(
        early_late_start_end_val_status5_cry_2_Y), .FCO(
        early_late_start_end_val_status5_cry_2_Z));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_14 (.A(
        early_found_msb_126_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[53]), .D(early_flags_msb_Z[117]), .FCI(
        early_found_msb_126_2_1_co0_6), .S(
        early_found_msb_126_2_1_wmux_14_S), .Y(
        early_found_msb_126_2_1_y3_0), .FCO(
        early_found_msb_126_2_1_co1_6));
    CFG3 #( .INIT(8'h08) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_i_a3_2_0[0]  (.A(
        clkalign_curr_state_Z[2]), .B(N_651), .C(N_523), .Y(
        wait_cnt_3_i_a3_2_0[0]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_40 (.A(
        late_found_msb_63_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[46]), .D(late_flags_msb_Z[110]), .FCI(
        late_found_msb_63_2_1_co0_19), .S(
        late_found_msb_63_2_1_wmux_40_S), .Y(
        late_found_msb_63_2_1_y5_2), .FCO(late_found_msb_63_2_1_co1_19)
        );
    SLE \late_flags_msb[81]  (.D(late_flags_msb_Z[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[81]));
    CFG2 #( .INIT(4'h2) )  
        \clkalign_curr_state_ns_5_0_.early_late_start_set5_0_a2  (.A(
        early_or_late_found_Z), .B(emflag_cnt_done_d_Z), .Y(N_653));
    CFG4 #( .INIT(16'h52EC) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_6_0_0_933_1  
        (.A(clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[3]), 
        .C(clkalign_curr_state_Z[1]), .D(clkalign_curr_state_Z[0]), .Y(
        un1_clkalign_curr_state_0_sqmuxa_6_0_0_933_1));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[8]), 
        .D(late_flags_msb_Z[72]), .FCI(late_found_msb_63_2_1_co1_0), 
        .S(late_found_msb_63_2_1_wmux_3_S), .Y(
        late_found_msb_63_2_1_y0_1), .FCO(late_found_msb_63_2_1_co0_1));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_21 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_63_2_1_co1_9), .S(
        early_found_msb_63_2_1_wmux_21_S), .Y(
        early_found_msb_63_2_1_wmux_21_Y), .FCO(
        early_found_msb_63_2_1_co0_10));
    SLE \early_flags_msb[78]  (.D(early_flags_msb_Z[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[78]));
    CFG4 #( .INIT(16'hCAC0) )  \clkalign_curr_state_ns_5_0_.m123  (.A(
        N_78), .B(N_118), .C(clkalign_curr_state_Z[5]), .D(m122_0_0), 
        .Y(clkalign_curr_state_ns[5]));
    CFG4 #( .INIT(16'h8CCC) )  
        \clkalign_curr_state_ns_5_0_.calc_done_0_sqmuxa_0_a3  (.A(
        emflag_cnt_done_d_Z), .B(clkalign_curr_state_d[27]), .C(
        N_538_i), .D(N_552_i), .Y(calc_done_0_sqmuxa));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_s[7]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[7]), .D(GND), .FCI(
        tap_cnt_cry_Z[6]), .S(tap_cnt_s_Z[7]), .Y(tap_cnt_s_Y[7]), 
        .FCO(tap_cnt_s_FCO[7]));
    SLE \late_flags_msb[35]  (.D(late_flags_msb_Z[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[35]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_30 (.A(
        early_found_lsb_63_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[58]), .D(early_flags_lsb_Z[122]), .FCI(
        early_found_lsb_63_2_1_co0_14), .S(
        early_found_lsb_63_2_1_wmux_30_S), .Y(
        early_found_lsb_63_2_1_y7_1), .FCO(
        early_found_lsb_63_2_1_co1_14));
    SLE \late_flags_lsb[37]  (.D(late_flags_lsb_Z[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[37]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_24 (.A(
        late_found_lsb_63_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[34]), .D(late_flags_lsb_Z[98]), .FCI(
        late_found_lsb_63_2_1_co0_11), .S(
        late_found_lsb_63_2_1_wmux_24_S), .Y(
        late_found_lsb_63_2_1_y1_1), .FCO(late_found_lsb_63_2_1_co1_11)
        );
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[7]), 
        .D(late_flags_lsb_Z[71]), .FCI(late_found_lsb_126_2_1_co1_16), 
        .S(late_found_lsb_126_2_1_wmux_35_S), .Y(
        late_found_lsb_126_2_1_y0_15), .FCO(
        late_found_lsb_126_2_1_co0_17));
    CFG4 #( .INIT(16'h3EED) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_o2_1_0[1]  (.A(
        clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[5]), .C(
        clkalign_curr_state_Z[4]), .D(clkalign_curr_state_Z[1]), .Y(
        N_537));
    CFG4 #( .INIT(16'hD1F3) )  \clkalign_curr_state_ns_5_0_.m92  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), .C(
        N_131_mux), .D(N_30), .Y(N_93));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[10])
        , .D(late_flags_lsb_Z[74]), .FCI(late_found_lsb_63_2_1_co1_12), 
        .S(late_found_lsb_63_2_1_wmux_27_S), .Y(
        late_found_lsb_63_2_1_y0_12), .FCO(
        late_found_lsb_63_2_1_co0_13));
    SLE \emflag_cnt[5]  (.D(emflag_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[5]));
    SLE \tapcnt_offset[1]  (.D(tapcnt_offset_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[1]));
    SLE \late_flags_lsb[44]  (.D(late_flags_lsb_Z[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[44]));
    SLE \tapcnt_offset[6]  (.D(tapcnt_offset_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[4])
        , .D(early_flags_msb_Z[68]), .FCI(early_found_msb_63_2_1_co1_4)
        , .S(early_found_msb_63_2_1_wmux_11_S), .Y(
        early_found_msb_63_2_1_y0_5), .FCO(
        early_found_msb_63_2_1_co0_5));
    SLE \early_flags_msb[69]  (.D(early_flags_msb_Z[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[69]));
    SLE \early_flags_msb[106]  (.D(early_flags_msb_Z[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[106]));
    SLE \early_late_init_val[7]  (.D(emflag_cnt_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[7]));
    SLE \tap_cnt[4]  (.D(tap_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[4]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_126_2_1_wmux_43 (.A(
        late_found_lsb_126_2_1_y7_2), .B(late_found_lsb_126_2_1_y5_2), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co1_20), .S(
        late_found_lsb_126_2_1_wmux_43_S), .Y(
        late_found_lsb_126_2_1_y0_19), .FCO(
        late_found_lsb_126_2_1_co0_21));
    SLE \late_flags_msb[85]  (.D(late_flags_msb_Z[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[85]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[7])
        , .D(early_flags_msb_Z[71]), .FCI(
        early_found_msb_126_2_1_co1_16), .S(
        early_found_msb_126_2_1_wmux_35_S), .Y(
        early_found_msb_126_2_1_y0_15), .FCO(
        early_found_msb_126_2_1_co0_17));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[5]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_6_S), 
        .Y(sig_tapcnt_final_1_3_Z[5]));
    SLE \early_flags_lsb[42]  (.D(early_flags_lsb_Z[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[42]));
    SLE \early_late_init_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[3]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_12 (.A(
        early_found_lsb_63_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[36]), .D(early_flags_lsb_Z[100]), .FCI(
        early_found_lsb_63_2_1_co0_5), .S(
        early_found_lsb_63_2_1_wmux_12_S), .Y(
        early_found_lsb_63_2_1_y1_0), .FCO(
        early_found_lsb_63_2_1_co1_5));
    SLE \late_flags_lsb[108]  (.D(late_flags_lsb_Z[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[108]));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_cry[5]  (.A(VCC), .B(
        timeout_cnt_Z[5]), .C(GND), .D(GND), .FCI(timeout_cnt_cry_Z[4])
        , .S(timeout_cnt_s[5]), .Y(timeout_cnt_cry_Y[5]), .FCO(
        timeout_cnt_cry_Z[5]));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNIKNK44[4]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[4]), 
        .D(GND), .FCI(tapcnt_offset_cry[3]), .S(tapcnt_offset_s[4]), 
        .Y(tapcnt_offset_RNIKNK44_Y[4]), .FCO(tapcnt_offset_cry[4]));
    SLE \tap_cnt[3]  (.D(tap_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[3]));
    SLE \late_flags_lsb[98]  (.D(late_flags_lsb_Z[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[98]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_4 
        (.A(early_late_end_val_Z[4]), .B(early_late_start_val_Z[4]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_3_Z), .S(
        early_late_start_end_val_status5_cry_4_S), .Y(
        early_late_start_end_val_status5_cry_4_Y), .FCO(
        early_late_start_end_val_status5_cry_4_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_63_2_1_wmux_7 (.A(
        early_found_msb_63_2_1_0_y7), .B(early_found_msb_63_2_1_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co1_2), .S(
        early_found_msb_63_2_1_wmux_7_S), .Y(
        early_found_msb_63_2_1_y0_3), .FCO(
        early_found_msb_63_2_1_co0_3));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[23]), .D(early_flags_lsb_Z[87]), .FCI(
        early_found_lsb_126_2_1_co1_17), .S(
        early_found_lsb_126_2_1_wmux_37_S), .Y(
        early_found_lsb_126_2_1_y0_16), .FCO(
        early_found_lsb_126_2_1_co0_18));
    SLE \timeout_cnt[2]  (.D(timeout_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[2]));
    SLE \late_flags_lsb[50]  (.D(late_flags_lsb_Z[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[50]));
    CFG2 #( .INIT(4'h8) )  no_early_and_late_found_msb (.A(
        early_not_found_msb_d_Z), .B(late_not_found_msb_d_Z), .Y(
        no_early_and_late_found_msb_Z));
    SLE \early_flags_msb[43]  (.D(early_flags_msb_Z[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[43]));
    SLE \early_flags_lsb[77]  (.D(early_flags_lsb_Z[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[77]));
    SLE \late_flags_lsb[22]  (.D(late_flags_lsb_Z[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[22]));
    SLE \late_flags_lsb[34]  (.D(late_flags_lsb_Z[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[34]));
    CFG2 #( .INIT(4'h8) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_17_0_a3_0  
        (.A(N_594_1), .B(rx_err_Z), .Y(N_594));
    ARI1 #( .INIT(20'h47700) )  \tap_cnt_cry_cy[0]  (.A(VCC), .B(
        clkalign_curr_state_Z[0]), .C(clkalign_curr_state_Z[2]), .D(
        GND), .FCI(VCC), .S(tap_cnt_cry_cy_S[0]), .Y(
        tap_cnt_cry_cy_Y[0]), .FCO(tap_cnt_cry_cy));
    SLE \late_flags_lsb[116]  (.D(late_flags_lsb_Z[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[116]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[3]), 
        .D(late_flags_lsb_Z[67]), .FCI(late_found_lsb_126_2_1_co1_10), 
        .S(late_found_lsb_126_2_1_wmux_23_S), .Y(
        late_found_lsb_126_2_1_y0_10), .FCO(
        late_found_lsb_126_2_1_co0_11));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_44 (.A(
        early_found_msb_63_2_1_y0_19), .B(early_found_msb_63_2_1_y3_2), 
        .C(early_found_msb_63_2_1_y1_2), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co0_21), .S(
        early_found_msb_63_2_1_wmux_44_S), .Y(
        early_found_msb_63_2_1_0_y45), .FCO(
        early_found_msb_63_2_1_co1_21));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[5]), 
        .D(late_flags_lsb_Z[69]), .FCI(late_found_lsb_126_2_1_co1_4), 
        .S(late_found_lsb_126_2_1_wmux_11_S), .Y(
        late_found_lsb_126_2_1_y0_5), .FCO(
        late_found_lsb_126_2_1_co0_5));
    SLE \late_flags_msb[91]  (.D(late_flags_msb_Z[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[91]));
    SLE \early_flags_msb[15]  (.D(early_flags_msb_Z[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[15]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_8 (.A(
        late_found_lsb_126_2_1_y0_3), .B(late_found_lsb_126_2_1_0_y3), 
        .C(late_found_lsb_126_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co0_3), .S(
        late_found_lsb_126_2_1_wmux_8_S), .Y(
        late_found_lsb_126_2_1_0_y9), .FCO(
        late_found_lsb_126_2_1_co1_3));
    SLE \rst_cnt[8]  (.D(rst_cnt_s[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[8]));
    SLE emflag_cnt_done_d (.D(emflag_cnt_done_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_done_d_Z));
    CFG4 #( .INIT(16'h0437) )  \clkalign_curr_state_ns_5_0_.m94  (.A(
        clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[5]), .C(
        N_93), .D(N_89), .Y(clkalign_curr_state_ns[2]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[4]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[4]), .D(early_late_init_val_Z[4]), .Y(
        tapcnt_final_11_iv_1[4]));
    SLE \late_flags_lsb[122]  (.D(late_flags_lsb_Z[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[122]));
    CFG3 #( .INIT(8'h08) )  
        \clkalign_curr_state_ns_5_0_.un1_RX_CLK_ALIGN_LOAD5_0_a3_1_1  
        (.A(clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[5]), 
        .C(clkalign_curr_state_Z[3]), .Y(
        un1_RX_CLK_ALIGN_LOAD5_0_a3_1_1));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[18])
        , .D(late_flags_lsb_Z[82]), .FCI(late_found_lsb_63_2_1_co1_11), 
        .S(late_found_lsb_63_2_1_wmux_25_S), .Y(
        late_found_lsb_63_2_1_y0_11), .FCO(
        late_found_lsb_63_2_1_co0_12));
    SLE \late_flags_msb[2]  (.D(late_flags_msb_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[2]));
    SLE \early_late_nxt_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[0]));
    SLE \late_flags_lsb[82]  (.D(late_flags_lsb_Z[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[82]));
    CFG4 #( .INIT(16'hDD1D) )  
        \clkalign_curr_state_ns_5_0_.m37_2_1_1_0  (.A(N_32_i), .B(
        current_state_0), .C(clkalign_curr_state_Z[4]), .D(N_4), .Y(
        m37_2_1_1_0));
    SLE \early_late_init_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[2]));
    SLE \early_late_init_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[5]));
    SLE \late_flags_msb[57]  (.D(late_flags_msb_Z[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[57]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_6 (.A(
        early_found_msb_63_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[56]), .D(early_flags_msb_Z[120]), .FCI(
        early_found_msb_63_2_1_co0_2), .S(
        early_found_msb_63_2_1_wmux_6_S), .Y(
        early_found_msb_63_2_1_0_y7), .FCO(
        early_found_msb_63_2_1_co1_2));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_28 (.A(
        early_found_lsb_63_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[42]), .D(early_flags_lsb_Z[106]), .FCI(
        early_found_lsb_63_2_1_co0_13), .S(
        early_found_lsb_63_2_1_wmux_28_S), .Y(
        early_found_lsb_63_2_1_y5_1), .FCO(
        early_found_lsb_63_2_1_co1_13));
    SLE \late_flags_msb[95]  (.D(late_flags_msb_Z[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[95]));
    ARI1 #( .INIT(20'h0CEC2) )  early_found_lsb_126_2_1_wmux_10 (.A(
        early_found_lsb_126_2_1_0_y21), .B(
        early_found_lsb_126_2_1_0_y9), .C(emflag_cnt_Z[2]), .D(
        emflag_cnt_Z[1]), .FCI(early_found_lsb_126_2_1_co0_4), .S(
        early_found_lsb_126_2_1_wmux_10_S), .Y(
        early_found_lsb_126_2_1_y0_4), .FCO(
        early_found_lsb_126_2_1_co1_4));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[14]), .D(early_flags_lsb_Z[78]), .FCI(
        early_found_lsb_63_2_1_co1_18), .S(
        early_found_lsb_63_2_1_wmux_39_S), .Y(
        early_found_lsb_63_2_1_y0_17), .FCO(
        early_found_lsb_63_2_1_co0_19));
    SLE \early_flags_lsb[6]  (.D(early_flags_lsb_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[6]));
    SLE \late_flags_lsb[11]  (.D(late_flags_lsb_Z[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[11]));
    SLE \early_flags_msb[118]  (.D(early_flags_msb_Z[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[118]));
    SLE \tap_cnt[2]  (.D(tap_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[2]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[11])
        , .D(late_flags_msb_Z[75]), .FCI(late_found_msb_126_2_1_co1_12)
        , .S(late_found_msb_126_2_1_wmux_27_S), .Y(
        late_found_msb_126_2_1_y0_12), .FCO(
        late_found_msb_126_2_1_co0_13));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_26 (.A(
        early_found_lsb_63_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[50]), .D(early_flags_lsb_Z[114]), .FCI(
        early_found_lsb_63_2_1_co0_12), .S(
        early_found_lsb_63_2_1_wmux_26_S), .Y(
        early_found_lsb_63_2_1_y3_1), .FCO(
        early_found_lsb_63_2_1_co1_12));
    SLE \early_flags_msb[93]  (.D(early_flags_msb_Z[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[93]));
    SLE \late_flags_msb[76]  (.D(late_flags_msb_Z[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[76]));
    SLE \late_flags_msb[62]  (.D(late_flags_msb_Z[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[62]));
    ARI1 #( .INIT(20'h0EA4A) )  early_found_lsb_126_2_1_wmux_9 (.A(
        early_found_lsb_126_2_1_0_y45), .B(
        early_found_lsb_126_2_1_y0_4), .C(
        early_found_lsb_126_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        early_found_lsb_126_2_1_co1_3), .S(
        early_found_lsb_126_2_1_wmux_9_S), .Y(N_1967), .FCO(
        early_found_lsb_126_2_1_co0_4));
    SLE \late_flags_msb[73]  (.D(late_flags_msb_Z[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[73]));
    SLE \late_flags_lsb[104]  (.D(late_flags_lsb_Z[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[104]));
    SLE \early_flags_msb[30]  (.D(early_flags_msb_Z[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[30]));
    SLE \late_flags_lsb[15]  (.D(late_flags_lsb_Z[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[15]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_36 (.A(
        early_found_lsb_126_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[39]), .D(early_flags_lsb_Z[103]), .FCI(
        early_found_lsb_126_2_1_co0_17), .S(
        early_found_lsb_126_2_1_wmux_36_S), .Y(
        early_found_lsb_126_2_1_y1_2), .FCO(
        early_found_lsb_126_2_1_co1_17));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[5]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[5]), .D(early_late_start_val_Z[5]), 
        .Y(tapcnt_final_11_iv_0[5]));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_7 (.A(
        early_late_end_val_Z[7]), .B(early_late_start_val_Z[7]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_6_Z), .S(
        un3_sig_tapcnt_final_1_cry_7_S), .Y(
        un3_sig_tapcnt_final_1_cry_7_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_7_Z));
    CFG2 #( .INIT(4'h8) )  \clkalign_curr_state_ns_5_0_.m44_0  (.A(
        N_30), .B(N_125_mux), .Y(m44_0));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_63_2_1_wmux_31 (.A(
        early_found_msb_63_2_1_y7_1), .B(early_found_msb_63_2_1_y5_1), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co1_14), .S(
        early_found_msb_63_2_1_wmux_31_S), .Y(
        early_found_msb_63_2_1_y0_14), .FCO(
        early_found_msb_63_2_1_co0_15));
    SLE early_late_init_and_nxt_set (.D(early_late_init_and_nxt_set5_Z)
        , .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_late_init_and_nxt_set_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[15]), .D(early_flags_lsb_Z[79]), .FCI(
        early_found_lsb_126_2_1_co1_18), .S(
        early_found_lsb_126_2_1_wmux_39_S), .Y(
        early_found_lsb_126_2_1_y0_17), .FCO(
        early_found_lsb_126_2_1_co0_19));
    SLE \early_flags_lsb[74]  (.D(early_flags_lsb_Z[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[74]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[6]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[6]), .D(early_late_init_val_Z[6]), .Y(
        tapcnt_final_11_iv_1[6]));
    SLE \early_flags_lsb[97]  (.D(early_flags_lsb_Z[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[97]));
    SLE \early_flags_lsb[45]  (.D(early_flags_lsb_Z[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[45]));
    SLE \late_flags_msb[54]  (.D(late_flags_msb_Z[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[54]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_12 (.A(
        late_found_msb_63_2_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[36]), .D(late_flags_msb_Z[100]), .FCI(
        late_found_msb_63_2_1_co0_5), .S(
        late_found_msb_63_2_1_wmux_12_S), .Y(
        late_found_msb_63_2_1_y1_0), .FCO(late_found_msb_63_2_1_co1_5));
    CFG2 #( .INIT(4'h8) )  \clkalign_curr_state_ns_5_0_.timeout_fg_3  
        (.A(timeout_cnt_Z[0]), .B(timeout_cnt_Z[1]), .Y(timeout_fg_3));
    SLE \late_flags_lsb[99]  (.D(late_flags_lsb_Z[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[99]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_18 (.A(
        early_found_lsb_63_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[60]), .D(early_flags_lsb_Z[124]), .FCI(
        early_found_lsb_63_2_1_co0_8), .S(
        early_found_lsb_63_2_1_wmux_18_S), .Y(
        early_found_lsb_63_2_1_y7_0), .FCO(
        early_found_lsb_63_2_1_co1_8));
    SLE \late_flags_lsb[103]  (.D(late_flags_lsb_Z[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[103]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[10]), .D(early_flags_lsb_Z[74]), .FCI(
        early_found_lsb_63_2_1_co1_12), .S(
        early_found_lsb_63_2_1_wmux_27_S), .Y(
        early_found_lsb_63_2_1_y0_12), .FCO(
        early_found_lsb_63_2_1_co0_13));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_0 (.A(
        late_found_lsb_126_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[33]), .D(late_flags_lsb_Z[97]), .FCI(
        late_found_lsb_126_2_1_0_co0), .S(
        late_found_lsb_126_2_1_wmux_0_S), .Y(
        late_found_lsb_126_2_1_0_y1), .FCO(
        late_found_lsb_126_2_1_0_co1));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_32 (.A(
        late_found_lsb_63_2_1_y0_14), .B(late_found_lsb_63_2_1_y3_1), 
        .C(late_found_lsb_63_2_1_y1_1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co0_15), .S(
        late_found_lsb_63_2_1_wmux_32_S), .Y(
        late_found_lsb_63_2_1_0_y33), .FCO(
        late_found_lsb_63_2_1_co1_15));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[7]), 
        .D(late_flags_msb_Z[71]), .FCI(late_found_msb_126_2_1_co1_16), 
        .S(late_found_msb_126_2_1_wmux_35_S), .Y(
        late_found_msb_126_2_1_y0_15), .FCO(
        late_found_msb_126_2_1_co0_17));
    SLE \late_flags_lsb[112]  (.D(late_flags_lsb_Z[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[112]));
    SLE \early_late_nxt_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[2]));
    SLE \early_flags_lsb[71]  (.D(early_flags_lsb_Z[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[71]));
    SLE \early_flags_msb[87]  (.D(early_flags_msb_Z[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[87]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_16 (.A(
        early_found_lsb_63_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[44]), .D(early_flags_lsb_Z[108]), .FCI(
        early_found_lsb_63_2_1_co0_7), .S(
        early_found_lsb_63_2_1_wmux_16_S), .Y(
        early_found_lsb_63_2_1_y5_0), .FCO(
        early_found_lsb_63_2_1_co1_7));
    CFG3 #( .INIT(8'hEC) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_15_0  (.A(
        early_late_start_set5_0_a3_1), .B(clkalign_curr_state_s9_0_a3), 
        .C(N_653), .Y(un1_clkalign_curr_state_15_0));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[3]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[3]), .D(early_late_start_val_Z[3]), 
        .Y(tapcnt_final_11_iv_0[3]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_44 (.A(
        early_found_lsb_126_2_1_y0_19), .B(
        early_found_lsb_126_2_1_y3_2), .C(early_found_lsb_126_2_1_y1_2)
        , .D(emflag_cnt_Z[3]), .FCI(early_found_lsb_126_2_1_co0_21), 
        .S(early_found_lsb_126_2_1_wmux_44_S), .Y(
        early_found_lsb_126_2_1_0_y45), .FCO(
        early_found_lsb_126_2_1_co1_21));
    CFG2 #( .INIT(4'h2) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s27_0_a2  (.A(
        N_634_i), .B(clkalign_curr_state_Z[0]), .Y(
        clkalign_curr_state_d[27]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_18 (.A(
        late_found_lsb_63_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[60]), .D(late_flags_lsb_Z[124]), .FCI(
        late_found_lsb_63_2_1_co0_8), .S(
        late_found_lsb_63_2_1_wmux_18_S), .Y(
        late_found_lsb_63_2_1_y7_0), .FCO(late_found_lsb_63_2_1_co1_8));
    SLE \early_flags_lsb[37]  (.D(early_flags_lsb_Z[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[37]));
    SLE \early_late_nxt_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[6]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_5 
        (.A(early_late_nxt_val_Z[5]), .B(early_late_init_val_Z[5]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_4_Z), 
        .S(early_late_init_nxt_val_status5_cry_5_S), .Y(
        early_late_init_nxt_val_status5_cry_5_Y), .FCO(
        early_late_init_nxt_val_status5_cry_5_Z));
    SLE \early_flags_msb[72]  (.D(early_flags_msb_Z[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[72]));
    SLE \early_flags_lsb[76]  (.D(early_flags_lsb_Z[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[76]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_20 (.A(
        late_found_lsb_63_2_1_y0_9), .B(late_found_lsb_63_2_1_y3_0), 
        .C(late_found_lsb_63_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co0_9), .S(
        late_found_lsb_63_2_1_wmux_20_S), .Y(
        late_found_lsb_63_2_1_0_y21), .FCO(late_found_lsb_63_2_1_co1_9)
        );
    SLE \early_flags_msb[27]  (.D(early_flags_msb_Z[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[27]));
    CFG3 #( .INIT(8'hB1) )  \clkalign_curr_state_ns_5_0_.m87  (.A(
        clkalign_curr_state_Z[2]), .B(N_83), .C(N_87), .Y(N_88));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_22 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_63_2_1_co0_10), .S(
        late_found_msb_63_2_1_wmux_22_S), .Y(
        late_found_msb_63_2_1_wmux_22_Y), .FCO(
        late_found_msb_63_2_1_co1_10));
    SLE \emflag_cnt[7]  (.D(emflag_cnt_s_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[7]));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[0]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_1_S), 
        .Y(sig_tapcnt_final_1_3_Z[0]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_20 (.A(
        early_found_msb_63_2_1_y0_9), .B(early_found_msb_63_2_1_y3_0), 
        .C(early_found_msb_63_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co0_9), .S(
        early_found_msb_63_2_1_wmux_20_S), .Y(
        early_found_msb_63_2_1_0_y21), .FCO(
        early_found_msb_63_2_1_co1_9));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[21])
        , .D(late_flags_lsb_Z[85]), .FCI(late_found_lsb_126_2_1_co1_5), 
        .S(late_found_lsb_126_2_1_wmux_13_S), .Y(
        late_found_lsb_126_2_1_y0_6), .FCO(
        late_found_lsb_126_2_1_co0_6));
    SLE \late_flags_msb[10]  (.D(late_flags_msb_Z[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[10]));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[5]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[5]), .D(GND), .FCI(
        tap_cnt_cry_Z[4]), .S(tap_cnt_s[5]), .Y(tap_cnt_cry_Y[5]), 
        .FCO(tap_cnt_cry_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[27])
        , .D(late_flags_lsb_Z[91]), .FCI(late_found_lsb_126_2_1_co1_13)
        , .S(late_found_lsb_126_2_1_wmux_29_S), .Y(
        late_found_lsb_126_2_1_y0_13), .FCO(
        late_found_lsb_126_2_1_co0_14));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_cry[2]  (.A(VCC), .B(
        timeout_cnt_Z[2]), .C(GND), .D(GND), .FCI(timeout_cnt_cry_Z[1])
        , .S(timeout_cnt_s[2]), .Y(timeout_cnt_cry_Y[2]), .FCO(
        timeout_cnt_cry_Z[2]));
    SLE \timeout_cnt[5]  (.D(timeout_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(timeout_cnt_Z[5]));
    SLE \emflag_cnt[1]  (.D(emflag_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[1]));
    SLE \late_flags_lsb[27]  (.D(late_flags_lsb_Z[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[27]));
    CFG3 #( .INIT(8'hE2) )  no_early_and_late_found (.A(
        no_early_and_late_found_lsb_d_Z), .B(emflag_cnt_Z[7]), .C(
        no_early_and_late_found_msb_d_Z), .Y(no_early_and_late_found_Z)
        );
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[28]), .D(early_flags_lsb_Z[92]), .FCI(
        early_found_lsb_63_2_1_co1_7), .S(
        early_found_lsb_63_2_1_wmux_17_S), .Y(
        early_found_lsb_63_2_1_y0_8), .FCO(
        early_found_lsb_63_2_1_co0_8));
    ARI1 #( .INIT(20'h0CEC2) )  early_found_msb_63_2_1_wmux_10 (.A(
        early_found_msb_63_2_1_0_y21), .B(early_found_msb_63_2_1_0_y9), 
        .C(emflag_cnt_Z[2]), .D(emflag_cnt_Z[1]), .FCI(
        early_found_msb_63_2_1_co0_4), .S(
        early_found_msb_63_2_1_wmux_10_S), .Y(
        early_found_msb_63_2_1_y0_4), .FCO(
        early_found_msb_63_2_1_co1_4));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_42 (.A(
        late_found_lsb_63_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[62]), .D(late_flags_lsb_Z[126]), .FCI(
        late_found_lsb_63_2_1_co0_20), .S(
        late_found_lsb_63_2_1_wmux_42_S), .Y(
        late_found_lsb_63_2_1_y7_2), .FCO(late_found_lsb_63_2_1_co1_20)
        );
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_14 (.A(
        late_found_msb_63_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[52]), .D(late_flags_msb_Z[116]), .FCI(
        late_found_msb_63_2_1_co0_6), .S(
        late_found_msb_63_2_1_wmux_14_S), .Y(
        late_found_msb_63_2_1_y3_0), .FCO(late_found_msb_63_2_1_co1_6));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[28])
        , .D(late_flags_msb_Z[92]), .FCI(late_found_msb_63_2_1_co1_7), 
        .S(late_found_msb_63_2_1_wmux_17_S), .Y(
        late_found_msb_63_2_1_y0_8), .FCO(late_found_msb_63_2_1_co0_8));
    SLE \late_flags_msb[22]  (.D(late_flags_msb_Z[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[22]));
    SLE \early_late_end_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[4]));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[5]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_6_S), 
        .Y(sig_tapcnt_final_2_3_Z[5]));
    ARI1 #( .INIT(20'h0EA4A) )  early_found_msb_63_2_1_wmux_9 (.A(
        early_found_msb_63_2_1_0_y45), .B(early_found_msb_63_2_1_y0_4), 
        .C(early_found_msb_63_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        early_found_msb_63_2_1_co1_3), .S(
        early_found_msb_63_2_1_wmux_9_S), .Y(N_2158), .FCO(
        early_found_msb_63_2_1_co0_4));
    SLE \late_flags_lsb[109]  (.D(late_flags_lsb_Z[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[109]));
    SLE \early_flags_msb[125]  (.D(early_flags_msb_Z[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[125]));
    SLE \early_flags_lsb[94]  (.D(early_flags_lsb_Z[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[94]));
    SLE \late_flags_lsb[41]  (.D(late_flags_lsb_Z[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[41]));
    SLE \early_flags_lsb[78]  (.D(early_flags_lsb_Z[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[78]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_34 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_63_2_1_co0_16), .S(
        late_found_lsb_63_2_1_wmux_34_S), .Y(
        late_found_lsb_63_2_1_wmux_34_Y), .FCO(
        late_found_lsb_63_2_1_co1_16));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[22])
        , .D(late_flags_lsb_Z[86]), .FCI(late_found_lsb_63_2_1_co1_17), 
        .S(late_found_lsb_63_2_1_wmux_37_S), .Y(
        late_found_lsb_63_2_1_y0_16), .FCO(
        late_found_lsb_63_2_1_co0_18));
    CFG2 #( .INIT(4'hE) )  early_or_late_found_msb (.A(
        early_found_msb_d_Z), .B(late_found_msb_d_Z), .Y(
        early_or_late_found_msb_Z));
    SLE \late_flags_lsb[87]  (.D(late_flags_lsb_Z[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[87]));
    CFG4 #( .INIT(16'h1000) )  sig_tapcnt_final_111 (.A(
        early_late_end_val_Z[1]), .B(early_late_end_val_Z[2]), .C(
        sig_tapcnt_final_111_4_Z), .D(sig_tapcnt_final_111_3_Z), .Y(
        sig_tapcnt_final_111_Z));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_32 (.A(
        late_found_msb_126_2_1_y0_14), .B(late_found_msb_126_2_1_y3_1), 
        .C(late_found_msb_126_2_1_y1_1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co0_15), .S(
        late_found_msb_126_2_1_wmux_32_S), .Y(
        late_found_msb_126_2_1_0_y33), .FCO(
        late_found_msb_126_2_1_co1_15));
    CFG1 #( .INIT(2'h1) )  \timeout_cnt_RNO[0]  (.A(timeout_cnt_Z[0]), 
        .Y(timeout_cnt_s[0]));
    SLE \early_flags_lsb[83]  (.D(early_flags_lsb_Z[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[83]));
    CFG4 #( .INIT(16'hFDF5) )  
        \clkalign_curr_state_ns_5_0_.tap_cnt9_i_RNIN6A01  (.A(N_490), 
        .B(clkalign_curr_state_Z[0]), .C(
        clkalign_curr_state_1_sqmuxa_1), .D(N_606_1), .Y(tap_cnte));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_38 (.A(
        late_found_msb_126_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[55]), .D(late_flags_msb_Z[119]), .FCI(
        late_found_msb_126_2_1_co0_18), .S(
        late_found_msb_126_2_1_wmux_38_S), .Y(
        late_found_msb_126_2_1_y3_2), .FCO(
        late_found_msb_126_2_1_co1_18));
    SLE \early_flags_msb[60]  (.D(early_flags_msb_Z[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[60]));
    SLE \late_flags_lsb[9]  (.D(late_flags_lsb_Z[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[9]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[27]), .D(early_flags_msb_Z[91]), .FCI(
        early_found_msb_126_2_1_co1_13), .S(
        early_found_msb_126_2_1_wmux_29_S), .Y(
        early_found_msb_126_2_1_y0_13), .FCO(
        early_found_msb_126_2_1_co0_14));
    SLE RX_RESET_LANE (.D(RX_RESET_LANE5), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_0_sqmuxa_3_0), .ALn(current_state_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[29])
        , .D(late_flags_msb_Z[93]), .FCI(late_found_msb_126_2_1_co1_7), 
        .S(late_found_msb_126_2_1_wmux_17_S), .Y(
        late_found_msb_126_2_1_y0_8), .FCO(
        late_found_msb_126_2_1_co0_8));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_38 (.A(
        early_found_lsb_126_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[55]), .D(early_flags_lsb_Z[119]), .FCI(
        early_found_lsb_126_2_1_co0_18), .S(
        early_found_lsb_126_2_1_wmux_38_S), .Y(
        early_found_lsb_126_2_1_y3_2), .FCO(
        early_found_lsb_126_2_1_co1_18));
    SLE \late_flags_lsb[45]  (.D(late_flags_lsb_Z[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[45]));
    SLE \early_flags_msb[84]  (.D(early_flags_msb_Z[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[84]));
    SLE \early_flags_lsb[91]  (.D(early_flags_lsb_Z[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[91]));
    CFG4 #( .INIT(16'hFEF1) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3[2]  (.A(wait_cnt_Z[1]), 
        .B(N_546), .C(N_540), .D(wait_cnt_Z[2]), .Y(wait_cnt_3[2]));
    SLE \early_flags_lsb[121]  (.D(early_flags_lsb_Z[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[121]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_4 (.A(
        early_found_lsb_63_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[40]), .D(early_flags_lsb_Z[104]), .FCI(
        early_found_lsb_63_2_1_co0_1), .S(
        early_found_lsb_63_2_1_wmux_4_S), .Y(
        early_found_lsb_63_2_1_0_y5), .FCO(
        early_found_lsb_63_2_1_co1_1));
    CFG3 #( .INIT(8'hB8) )  \clkalign_curr_state_ns_5_0_.m88  (.A(N_88)
        , .B(clkalign_curr_state_Z[3]), .C(N_143_mux), .Y(N_89));
    CFG4 #( .INIT(16'h7BDE) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state63_NE_0  (.A(
        tapcnt_final_Z[6]), .B(tapcnt_final_Z[5]), .C(tap_cnt_Z[6]), 
        .D(tap_cnt_Z[5]), .Y(clkalign_curr_state63_NE_0));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_24 (.A(
        late_found_msb_63_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[34]), .D(late_flags_msb_Z[98]), .FCI(
        late_found_msb_63_2_1_co0_11), .S(
        late_found_msb_63_2_1_wmux_24_S), .Y(
        late_found_msb_63_2_1_y1_1), .FCO(late_found_msb_63_2_1_co1_11)
        );
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_38 (.A(
        late_found_lsb_126_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[55]), .D(late_flags_lsb_Z[119]), .FCI(
        late_found_lsb_126_2_1_co0_18), .S(
        late_found_lsb_126_2_1_wmux_38_S), .Y(
        late_found_lsb_126_2_1_y3_2), .FCO(
        late_found_lsb_126_2_1_co1_18));
    CFG4 #( .INIT(16'h8000) )  
        \clkalign_curr_state_ns_5_0_.timeout_fg  (.A(timeout_cnt_Z[3]), 
        .B(timeout_cnt_Z[2]), .C(timeout_fg_4), .D(timeout_fg_3), .Y(
        timeout_fg));
    CFG4 #( .INIT(16'h8000) )  
        \clkalign_curr_state_ns_5_0_.reset_dly_fg4_6  (.A(rst_cnt_Z[5])
        , .B(rst_cnt_Z[4]), .C(rst_cnt_Z[3]), .D(rst_cnt_Z[2]), .Y(
        reset_dly_fg4_6));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[10])
        , .D(late_flags_msb_Z[74]), .FCI(late_found_msb_63_2_1_co1_12), 
        .S(late_found_msb_63_2_1_wmux_27_S), .Y(
        late_found_msb_63_2_1_y0_12), .FCO(
        late_found_msb_63_2_1_co0_13));
    SLE \late_flags_lsb[24]  (.D(late_flags_lsb_Z[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[24]));
    SLE \early_flags_lsb[34]  (.D(early_flags_lsb_Z[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[34]));
    SLE \early_flags_msb[105]  (.D(early_flags_msb_Z[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[105]));
    SLE RX_CLK_ALIGN_ERR (.D(timeout_fg), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(CLK_TRAIN_ERROR_c));
    ARI1 #( .INIT(20'h4AA00) )  timeout_cnt_s_1134 (.A(VCC), .B(
        timeout_cnt_Z[0]), .C(GND), .D(GND), .FCI(VCC), .S(
        timeout_cnt_s_1134_S), .Y(timeout_cnt_s_1134_Y), .FCO(
        timeout_cnt_s_1134_FCO));
    SLE \late_flags_msb[67]  (.D(late_flags_msb_Z[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[67]));
    CFG4 #( .INIT(16'h3928) )  \clkalign_curr_state_ns_5_0_.m74  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), .C(
        m74_1_0), .D(N_32_i), .Y(N_75));
    SLE \early_flags_lsb[96]  (.D(early_flags_lsb_Z[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[96]));
    SLE \early_flags_msb[24]  (.D(early_flags_msb_Z[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[24]));
    SLE \late_flags_lsb[31]  (.D(late_flags_lsb_Z[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[31]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_24 (.A(
        early_found_lsb_126_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[35]), .D(early_flags_lsb_Z[99]), .FCI(
        early_found_lsb_126_2_1_co0_11), .S(
        early_found_lsb_126_2_1_wmux_24_S), .Y(
        early_found_lsb_126_2_1_y1_1), .FCO(
        early_found_lsb_126_2_1_co1_11));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[16])
        , .D(late_flags_lsb_Z[80]), .FCI(late_found_lsb_63_2_1_0_co1), 
        .S(late_found_lsb_63_2_1_wmux_1_S), .Y(
        late_found_lsb_63_2_1_y0_0), .FCO(late_found_lsb_63_2_1_co0_0));
    SLE \early_flags_msb[81]  (.D(early_flags_msb_Z[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[81]));
    SLE \early_flags_msb[120]  (.D(early_flags_msb_Z[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[120]));
    CFG2 #( .INIT(4'h8) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0_1  
        (.A(N_656), .B(N_639), .Y(
        un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0));
    SLE \sig_tapcnt_final_2[4]  (.D(sig_tapcnt_final_2_3_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[4]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_44 (.A(
        late_found_lsb_63_2_1_y0_19), .B(late_found_lsb_63_2_1_y3_2), 
        .C(late_found_lsb_63_2_1_y1_2), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co0_21), .S(
        late_found_lsb_63_2_1_wmux_44_S), .Y(
        late_found_lsb_63_2_1_0_y45), .FCO(
        late_found_lsb_63_2_1_co1_21));
    SLE \early_late_nxt_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[5]));
    CFG2 #( .INIT(4'h8) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s25_0_a2  (.A(
        clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[2]), .Y(
        N_639));
    SLE \late_flags_lsb[84]  (.D(late_flags_lsb_Z[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[84]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_34 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_63_2_1_co0_16), .S(
        early_found_lsb_63_2_1_wmux_34_S), .Y(
        early_found_lsb_63_2_1_wmux_34_Y), .FCO(
        early_found_lsb_63_2_1_co1_16));
    CFG4 #( .INIT(16'h8000) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_8_0_a2  
        (.A(N_2979), .B(N_627), .C(CO0_0), .D(cnt_Z[1]), .Y(N_643));
    CFG4 #( .INIT(16'h158C) )  \clkalign_curr_state_ns_5_0_.m104_1_2  
        (.A(clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), 
        .C(N_102), .D(N_82_i), .Y(m104_1_2));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[12])
        , .D(late_flags_msb_Z[76]), .FCI(late_found_msb_63_2_1_co1_6), 
        .S(late_found_msb_63_2_1_wmux_15_S), .Y(
        late_found_msb_63_2_1_y0_7), .FCO(late_found_msb_63_2_1_co0_7));
    SLE \late_flags_lsb[100]  (.D(late_flags_lsb_Z[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[100]));
    SLE \early_flags_lsb[69]  (.D(early_flags_lsb_Z[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[69]));
    SLE \early_flags_lsb[31]  (.D(early_flags_lsb_Z[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[31]));
    CFG3 #( .INIT(8'h08) )  
        \clkalign_curr_state_ns_5_0_.un1_RX_CLK_ALIGN_LOAD5_0_a3_1  (
        .A(N_642), .B(un1_RX_CLK_ALIGN_LOAD5_0_a3_1_1), .C(N_525), .Y(
        N_607));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_4 (.A(
        early_found_msb_126_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[41]), .D(early_flags_msb_Z[105]), .FCI(
        early_found_msb_126_2_1_co0_1), .S(
        early_found_msb_126_2_1_wmux_4_S), .Y(
        early_found_msb_126_2_1_0_y5), .FCO(
        early_found_msb_126_2_1_co1_1));
    SLE \early_flags_lsb[101]  (.D(early_flags_lsb_Z[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[101]));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[4]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_5_S), 
        .Y(sig_tapcnt_final_2_3_Z[4]));
    SLE \late_flags_msb[102]  (.D(late_flags_msb_Z[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[102]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[26]), .D(early_flags_msb_Z[90]), .FCI(
        early_found_msb_63_2_1_co1_13), .S(
        early_found_msb_63_2_1_wmux_29_S), .Y(
        early_found_msb_63_2_1_y0_13), .FCO(
        early_found_msb_63_2_1_co0_14));
    SLE \early_flags_msb[75]  (.D(early_flags_msb_Z[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[75]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_4 (.A(
        late_found_msb_63_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[40]), .D(late_flags_msb_Z[104]), .FCI(
        late_found_msb_63_2_1_co0_1), .S(
        late_found_msb_63_2_1_wmux_4_S), .Y(late_found_msb_63_2_1_0_y5)
        , .FCO(late_found_msb_63_2_1_co1_1));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_4 (.A(
        late_found_msb_126_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[41]), .D(late_flags_msb_Z[105]), .FCI(
        late_found_msb_126_2_1_co0_1), .S(
        late_found_msb_126_2_1_wmux_4_S), .Y(
        late_found_msb_126_2_1_0_y5), .FCO(
        late_found_msb_126_2_1_co1_1));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_16 (.A(
        early_found_msb_126_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[45]), .D(early_flags_msb_Z[109]), .FCI(
        early_found_msb_126_2_1_co0_7), .S(
        early_found_msb_126_2_1_wmux_16_S), .Y(
        early_found_msb_126_2_1_y5_0), .FCO(
        early_found_msb_126_2_1_co1_7));
    SLE \early_flags_msb[86]  (.D(early_flags_msb_Z[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[86]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[6]), 
        .D(late_flags_lsb_Z[70]), .FCI(late_found_lsb_63_2_1_co1_16), 
        .S(late_found_lsb_63_2_1_wmux_35_S), .Y(
        late_found_lsb_63_2_1_y0_15), .FCO(
        late_found_lsb_63_2_1_co0_17));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[9])
        , .D(early_flags_lsb_Z[73]), .FCI(
        early_found_lsb_126_2_1_co1_0), .S(
        early_found_lsb_126_2_1_wmux_3_S), .Y(
        early_found_lsb_126_2_1_y0_1), .FCO(
        early_found_lsb_126_2_1_co0_1));
    SLE \early_flags_msb[21]  (.D(early_flags_msb_Z[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[21]));
    SLE \early_flags_lsb[116]  (.D(early_flags_lsb_Z[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[116]));
    SLE \late_flags_lsb[35]  (.D(late_flags_lsb_Z[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[35]));
    ARI1 #( .INIT(20'h0EA4A) )  late_found_msb_63_2_1_wmux_9 (.A(
        late_found_msb_63_2_1_0_y45), .B(late_found_msb_63_2_1_y0_4), 
        .C(late_found_msb_63_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        late_found_msb_63_2_1_co1_3), .S(
        late_found_msb_63_2_1_wmux_9_S), .Y(N_2285), .FCO(
        late_found_msb_63_2_1_co0_4));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[25])
        , .D(late_flags_lsb_Z[89]), .FCI(late_found_lsb_126_2_1_co1_1), 
        .S(late_found_lsb_126_2_1_wmux_5_S), .Y(
        late_found_lsb_126_2_1_y0_2), .FCO(
        late_found_lsb_126_2_1_co0_2));
    CFG2 #( .INIT(4'h8) )  early_late_init_and_nxt_set5 (.A(
        early_late_init_set_Z), .B(early_late_nxt_set_Z), .Y(
        early_late_init_and_nxt_set5_Z));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_8 (.A(
        late_found_lsb_63_2_1_y0_3), .B(late_found_lsb_63_2_1_0_y3), 
        .C(late_found_lsb_63_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co0_3), .S(
        late_found_lsb_63_2_1_wmux_8_S), .Y(late_found_lsb_63_2_1_0_y9)
        , .FCO(late_found_lsb_63_2_1_co1_3));
    SLE \late_flags_msb[126]  (.D(late_flags_msb_Z[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[126]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[6]  (.A(VCC), .B(
        rst_cnt_Z[6]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[5]), .S(
        rst_cnt_s[6]), .Y(rst_cnt_cry_Y[6]), .FCO(rst_cnt_cry_Z[6]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_63_2_1_wmux_19 (.A(
        early_found_msb_63_2_1_y7_0), .B(early_found_msb_63_2_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_63_2_1_co1_8), .S(
        early_found_msb_63_2_1_wmux_19_S), .Y(
        early_found_msb_63_2_1_y0_9), .FCO(
        early_found_msb_63_2_1_co0_9));
    SLE \early_flags_lsb[36]  (.D(early_flags_lsb_Z[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[36]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_126_2_1_wmux_31 (.A(
        early_found_msb_126_2_1_y7_1), .B(early_found_msb_126_2_1_y5_1)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_126_2_1_co1_14), .S(
        early_found_msb_126_2_1_wmux_31_S), .Y(
        early_found_msb_126_2_1_y0_14), .FCO(
        early_found_msb_126_2_1_co0_15));
    SLE \early_flags_lsb[98]  (.D(early_flags_lsb_Z[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[98]));
    CFG3 #( .INIT(8'h08) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_11_0_a2  
        (.A(clkalign_curr_state_Z[2]), .B(N_627), .C(N_523), .Y(
        N_634_i));
    CFG4 #( .INIT(16'h8000) )  
        \clkalign_curr_state_ns_5_0_.timeout_fg_4  (.A(
        timeout_cnt_Z[7]), .B(timeout_cnt_Z[6]), .C(timeout_cnt_Z[5]), 
        .D(timeout_cnt_Z[4]), .Y(timeout_fg_4));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_44 (.A(
        late_found_msb_126_2_1_y0_19), .B(late_found_msb_126_2_1_y3_2), 
        .C(late_found_msb_126_2_1_y1_2), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co0_21), .S(
        late_found_msb_126_2_1_wmux_44_S), .Y(
        late_found_msb_126_2_1_0_y45), .FCO(
        late_found_msb_126_2_1_co1_21));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_63_2_1_wmux_7 (.A(
        late_found_lsb_63_2_1_0_y7), .B(late_found_lsb_63_2_1_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_63_2_1_co1_2), .S(
        late_found_lsb_63_2_1_wmux_7_S), .Y(late_found_lsb_63_2_1_y0_3)
        , .FCO(late_found_lsb_63_2_1_co0_3));
    CFG3 #( .INIT(8'hB1) )  \clkalign_curr_state_ns_5_0_.m118  (.A(
        clkalign_curr_state_Z[5]), .B(N_116), .C(N_118), .Y(
        clkalign_curr_state_ns[4]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_40 (.A(
        late_found_lsb_126_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[47]), .D(late_flags_lsb_Z[111]), .FCI(
        late_found_lsb_126_2_1_co0_19), .S(
        late_found_lsb_126_2_1_wmux_40_S), .Y(
        late_found_lsb_126_2_1_y5_2), .FCO(
        late_found_lsb_126_2_1_co1_19));
    CFG3 #( .INIT(8'hEC) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_end_set12_1_0  (.A(
        un1_early_late_end_set12_1_0_a3_1), .B(
        clkalign_curr_state_s9_0_a3), .C(N_653), .Y(
        un1_early_late_end_set12_1_0));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_4 (.A(
        early_late_end_val_Z[4]), .B(early_late_start_val_Z[4]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_3_Z), .S(
        un3_sig_tapcnt_final_1_cry_4_S), .Y(
        un3_sig_tapcnt_final_1_cry_4_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_4_Z));
    SLE \early_flags_msb[26]  (.D(early_flags_msb_Z[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[26]));
    SLE \early_flags_msb[100]  (.D(early_flags_msb_Z[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[100]));
    SLE \early_flags_lsb[29]  (.D(early_flags_lsb_Z[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[29]));
    CFG4 #( .INIT(16'h8000) )  \clkalign_curr_state_ns_5_0_.m86_3  (.A(
        clkalign_curr_state_Z[4]), .B(N_60), .C(
        no_early_and_late_found_Z), .D(clkalign_curr_state_Z[1]), .Y(
        m86_2));
    SLE \late_flags_msb[64]  (.D(late_flags_msb_Z[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[64]));
    SLE \sig_tapcnt_final_2[6]  (.D(sig_tapcnt_final_2_3_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[6]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_6 (.A(
        late_found_lsb_63_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[56]), .D(late_flags_lsb_Z[120]), .FCI(
        late_found_lsb_63_2_1_co0_2), .S(
        late_found_lsb_63_2_1_wmux_6_S), .Y(late_found_lsb_63_2_1_0_y7)
        , .FCO(late_found_lsb_63_2_1_co1_2));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_6 (.A(
        early_found_msb_126_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[57]), .D(early_flags_msb_Z[121]), .FCI(
        early_found_msb_126_2_1_co0_2), .S(
        early_found_msb_126_2_1_wmux_6_S), .Y(
        early_found_msb_126_2_1_0_y7), .FCO(
        early_found_msb_126_2_1_co1_2));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[18])
        , .D(late_flags_msb_Z[82]), .FCI(late_found_msb_63_2_1_co1_11), 
        .S(late_found_msb_63_2_1_wmux_25_S), .Y(
        late_found_msb_63_2_1_y0_11), .FCO(
        late_found_msb_63_2_1_co0_12));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_30 (.A(
        early_found_msb_63_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[58]), .D(early_flags_msb_Z[122]), .FCI(
        early_found_msb_63_2_1_co0_14), .S(
        early_found_msb_63_2_1_wmux_30_S), .Y(
        early_found_msb_63_2_1_y7_1), .FCO(
        early_found_msb_63_2_1_co1_14));
    SLE \late_flags_msb[8]  (.D(late_flags_msb_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[8]));
    SLE \emflag_cnt[0]  (.D(emflag_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[0]));
    SLE \late_flags_lsb[58]  (.D(late_flags_lsb_Z[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[58]));
    SLE \early_flags_msb[88]  (.D(early_flags_msb_Z[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[88]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_126_2_1_wmux_19 (.A(
        late_found_lsb_126_2_1_y7_0), .B(late_found_lsb_126_2_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co1_8), .S(
        late_found_lsb_126_2_1_wmux_19_S), .Y(
        late_found_lsb_126_2_1_y0_9), .FCO(
        late_found_lsb_126_2_1_co0_9));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_2 (.A(
        late_found_msb_126_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[49]), .D(late_flags_msb_Z[113]), .FCI(
        late_found_msb_126_2_1_co0_0), .S(
        late_found_msb_126_2_1_wmux_2_S), .Y(
        late_found_msb_126_2_1_0_y3), .FCO(
        late_found_msb_126_2_1_co1_0));
    SLE \early_flags_lsb[38]  (.D(early_flags_lsb_Z[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[38]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_126_2_1_wmux_43 (.A(
        early_found_lsb_126_2_1_y7_2), .B(early_found_lsb_126_2_1_y5_2)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_126_2_1_co1_20), .S(
        early_found_lsb_126_2_1_wmux_43_S), .Y(
        early_found_lsb_126_2_1_y0_19), .FCO(
        early_found_lsb_126_2_1_co0_21));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[24]), .D(early_flags_msb_Z[88]), .FCI(
        early_found_msb_63_2_1_co1_1), .S(
        early_found_msb_63_2_1_wmux_5_S), .Y(
        early_found_msb_63_2_1_y0_2), .FCO(
        early_found_msb_63_2_1_co0_2));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_24 (.A(
        late_found_msb_126_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[35]), .D(late_flags_msb_Z[99]), .FCI(
        late_found_msb_126_2_1_co0_11), .S(
        late_found_msb_126_2_1_wmux_24_S), .Y(
        late_found_msb_126_2_1_y1_1), .FCO(
        late_found_msb_126_2_1_co1_11));
    SLE \late_flags_msb[70]  (.D(late_flags_msb_Z[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[70]));
    SLE \early_flags_msb[28]  (.D(early_flags_msb_Z[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[28]));
    SLE \late_flags_msb[51]  (.D(late_flags_msb_Z[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[51]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_20 (.A(
        late_found_lsb_126_2_1_y0_9), .B(late_found_lsb_126_2_1_y3_0), 
        .C(late_found_lsb_126_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co0_9), .S(
        late_found_lsb_126_2_1_wmux_20_S), .Y(
        late_found_lsb_126_2_1_0_y21), .FCO(
        late_found_lsb_126_2_1_co1_9));
    SLE \late_flags_lsb[6]  (.D(late_flags_lsb_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[6]));
    SLE \late_flags_msb[6]  (.D(late_flags_msb_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[6]));
    CFG4 #( .INIT(16'h0200) )  
        \clkalign_curr_state_ns_5_0_.timeout_cnt10_0_a3  (.A(
        clkalign_curr_state_d[27]), .B(early_late_init_and_nxt_set_Z), 
        .C(early_late_start_and_end_set_Z), .D(emflag_cnt_done_d_Z), 
        .Y(timeout_cnte));
    SLE \late_flags_msb[27]  (.D(late_flags_msb_Z[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[27]));
    SLE \late_flags_lsb[72]  (.D(late_flags_lsb_Z[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[72]));
    SLE \late_flags_msb[118]  (.D(late_flags_msb_Z[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[118]));
    SLE \late_flags_msb[9]  (.D(late_flags_msb_Z[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[9]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_26 (.A(
        late_found_msb_126_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[51]), .D(late_flags_msb_Z[115]), .FCI(
        late_found_msb_126_2_1_co0_12), .S(
        late_found_msb_126_2_1_wmux_26_S), .Y(
        late_found_msb_126_2_1_y3_1), .FCO(
        late_found_msb_126_2_1_co1_12));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[3]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[3]), .D(early_late_init_val_Z[3]), .Y(
        tapcnt_final_11_iv_1[3]));
    SLE \rst_cnt[7]  (.D(rst_cnt_s[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[7]));
    CFG4 #( .INIT(16'h0400) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_8_0_a3_0  
        (.A(N_525), .B(N_125_mux), .C(clkalign_curr_state_Z[5]), .D(
        N_2979), .Y(N_622));
    CFG4 #( .INIT(16'hBCB0) )  \clkalign_curr_state_ns_5_0_.m16_2  (.A(
        N_5), .B(clkalign_curr_state_Z[1]), .C(m16_1), .D(N_4), .Y(
        m16_2));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[31]), .D(early_flags_lsb_Z[95]), .FCI(
        early_found_lsb_126_2_1_co1_19), .S(
        early_found_lsb_126_2_1_wmux_41_S), .Y(
        early_found_lsb_126_2_1_y0_18), .FCO(
        early_found_lsb_126_2_1_co0_20));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_0 (.A(
        early_found_lsb_126_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[33]), .D(early_flags_lsb_Z[97]), .FCI(
        early_found_lsb_126_2_1_0_co0), .S(
        early_found_lsb_126_2_1_wmux_0_S), .Y(
        early_found_lsb_126_2_1_0_y1), .FCO(
        early_found_lsb_126_2_1_0_co1));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_cry[6]  (.A(VCC), .B(
        timeout_cnt_Z[6]), .C(GND), .D(GND), .FCI(timeout_cnt_cry_Z[5])
        , .S(timeout_cnt_s[6]), .Y(timeout_cnt_cry_Y[6]), .FCO(
        timeout_cnt_cry_Z[6]));
    SLE \late_flags_msb[55]  (.D(late_flags_msb_Z[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[55]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_126_2_1_wmux_31 (.A(
        late_found_lsb_126_2_1_y7_1), .B(late_found_lsb_126_2_1_y5_1), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co1_14), .S(
        late_found_lsb_126_2_1_wmux_31_S), .Y(
        late_found_lsb_126_2_1_y0_14), .FCO(
        late_found_lsb_126_2_1_co0_15));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_8 (.A(
        early_found_msb_126_2_1_y0_3), .B(early_found_msb_126_2_1_0_y3)
        , .C(early_found_msb_126_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_126_2_1_co0_3), .S(
        early_found_msb_126_2_1_wmux_8_S), .Y(
        early_found_msb_126_2_1_0_y9), .FCO(
        early_found_msb_126_2_1_co1_3));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_2 (.A(
        early_found_msb_126_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[49]), .D(early_flags_msb_Z[113]), .FCI(
        early_found_msb_126_2_1_co0_0), .S(
        early_found_msb_126_2_1_wmux_2_S), .Y(
        early_found_msb_126_2_1_0_y3), .FCO(
        early_found_msb_126_2_1_co1_0));
    CFG2 #( .INIT(4'hD) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_1_sqmuxa_2_0_o2  
        (.A(early_late_start_and_end_set_Z), .B(
        tapcnt_final_1_status_Z), .Y(N_538_i));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[2]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_3_S), 
        .Y(sig_tapcnt_final_1_3_Z[2]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_28 (.A(
        late_found_lsb_63_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[42]), .D(late_flags_lsb_Z[106]), .FCI(
        late_found_lsb_63_2_1_co0_13), .S(
        late_found_lsb_63_2_1_wmux_28_S), .Y(
        late_found_lsb_63_2_1_y5_1), .FCO(late_found_lsb_63_2_1_co1_13)
        );
    SLE \late_flags_msb[116]  (.D(late_flags_msb_Z[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[116]));
    CFG2 #( .INIT(4'h2) )  \clkalign_curr_state_ns_5_0_.m29  (.A(
        clkalign_curr_state_Z[4]), .B(clkalign_curr_state_Z[0]), .Y(
        N_30));
    SLE RX_CLK_ALIGN_MOVE (.D(N_2924_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_1_sqmuxa_5_0), .ALn(current_state_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV));
    ARI1 #( .INIT(20'h0CEC2) )  late_found_msb_63_2_1_wmux_10 (.A(
        late_found_msb_63_2_1_0_y21), .B(late_found_msb_63_2_1_0_y9), 
        .C(emflag_cnt_Z[2]), .D(emflag_cnt_Z[1]), .FCI(
        late_found_msb_63_2_1_co0_4), .S(
        late_found_msb_63_2_1_wmux_10_S), .Y(
        late_found_msb_63_2_1_y0_4), .FCO(late_found_msb_63_2_1_co1_4));
    SLE \early_flags_msb[59]  (.D(early_flags_msb_Z[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[59]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_30 (.A(
        late_found_lsb_63_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[58]), .D(late_flags_lsb_Z[122]), .FCI(
        late_found_lsb_63_2_1_co0_14), .S(
        late_found_lsb_63_2_1_wmux_30_S), .Y(
        late_found_lsb_63_2_1_y7_1), .FCO(late_found_lsb_63_2_1_co1_14)
        );
    SLE \early_flags_lsb[72]  (.D(early_flags_lsb_Z[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[72]));
    CFG2 #( .INIT(4'hE) )  clkalign_curr_state81_NE_3 (.A(
        tapcnt_offset_Z[6]), .B(tapcnt_offset_Z[7]), .Y(
        clkalign_curr_state81_NE_3_Z));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[0]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_1_S), 
        .Y(sig_tapcnt_final_2_3_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_40 (.A(
        early_found_msb_126_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[47]), .D(early_flags_msb_Z[111]), .FCI(
        early_found_msb_126_2_1_co0_19), .S(
        early_found_msb_126_2_1_wmux_40_S), .Y(
        early_found_msb_126_2_1_y5_2), .FCO(
        early_found_msb_126_2_1_co1_19));
    SLE rx_err (.D(timeout_cnte), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(un1_clkalign_curr_state_17_0), .ALn(current_state_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_err_Z));
    SLE \late_flags_msb[24]  (.D(late_flags_msb_Z[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[24]));
    SLE \early_flags_msb[8]  (.D(early_flags_msb_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[8]));
    CFG1 #( .INIT(2'h1) )  \cnt_RNO[0]  (.A(CO0_0), .Y(CO0_0_i));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[13]), .D(early_flags_msb_Z[77]), .FCI(
        early_found_msb_126_2_1_co1_6), .S(
        early_found_msb_126_2_1_wmux_15_S), .Y(
        early_found_msb_126_2_1_y0_7), .FCO(
        early_found_msb_126_2_1_co0_7));
    SLE \early_flags_lsb[110]  (.D(early_flags_lsb_Z[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[110]));
    SLE \rst_cnt[0]  (.D(rst_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[14]), .D(early_flags_msb_Z[78]), .FCI(
        early_found_msb_63_2_1_co1_18), .S(
        early_found_msb_63_2_1_wmux_39_S), .Y(
        early_found_msb_63_2_1_y0_17), .FCO(
        early_found_msb_63_2_1_co0_19));
    SLE \early_flags_msb[37]  (.D(early_flags_msb_Z[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[37]));
    CFG4 #( .INIT(16'hCCEC) )  
        \clkalign_curr_state_ns_5_0_.RX_RESET_LANE5_0_o3  (.A(N_656), 
        .B(N_585_i), .C(clkalign_curr_state_Z[2]), .D(N_523), .Y(
        RX_RESET_LANE5));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_20 (.A(
        late_found_msb_63_2_1_y0_9), .B(late_found_msb_63_2_1_y3_0), 
        .C(late_found_msb_63_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co0_9), .S(
        late_found_msb_63_2_1_wmux_20_S), .Y(
        late_found_msb_63_2_1_0_y21), .FCO(late_found_msb_63_2_1_co1_9)
        );
    SLE \early_flags_lsb[13]  (.D(early_flags_lsb_Z[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[13]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[29]), .D(early_flags_lsb_Z[93]), .FCI(
        early_found_lsb_126_2_1_co1_7), .S(
        early_found_lsb_126_2_1_wmux_17_S), .Y(
        early_found_lsb_126_2_1_y0_8), .FCO(
        early_found_lsb_126_2_1_co0_8));
    CFG4 #( .INIT(16'hFFF8) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_0_sqmuxa_4_0_a3_0_RNIRB5O  
        (.A(clkalign_curr_state_0_sqmuxa_4_0_a3_0), .B(N_642), .C(
        clkalign_curr_state_s9_0_a3), .D(clkalign_curr_state_d[27]), 
        .Y(tapcnt_offsete));
    SLE \late_flags_lsb[59]  (.D(late_flags_lsb_Z[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[59]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_4 (.A(
        early_found_msb_63_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[40]), .D(early_flags_msb_Z[104]), .FCI(
        early_found_msb_63_2_1_co0_1), .S(
        early_found_msb_63_2_1_wmux_4_S), .Y(
        early_found_msb_63_2_1_0_y5), .FCO(
        early_found_msb_63_2_1_co1_1));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[3])
        , .D(early_flags_lsb_Z[67]), .FCI(
        early_found_lsb_126_2_1_co1_10), .S(
        early_found_lsb_126_2_1_wmux_23_S), .Y(
        early_found_lsb_126_2_1_y0_10), .FCO(
        early_found_lsb_126_2_1_co0_11));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[6]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[6]), .D(GND), .FCI(
        tap_cnt_cry_Z[5]), .S(tap_cnt_s[6]), .Y(tap_cnt_cry_Y[6]), 
        .FCO(tap_cnt_cry_Z[6]));
    CFG4 #( .INIT(16'hB975) )  \clkalign_curr_state_ns_5_0_.m57  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[4]), .C(
        N_19_i), .D(m57_1_2), .Y(N_58));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[4]  (.A(VCC), .B(
        rst_cnt_Z[4]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[3]), .S(
        rst_cnt_s[4]), .Y(rst_cnt_cry_Y[4]), .FCO(rst_cnt_cry_Z[4]));
    SLE \late_flags_lsb[4]  (.D(late_flags_lsb_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[4]));
    SLE \early_flags_msb[112]  (.D(early_flags_msb_Z[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[112]));
    SLE \early_flags_lsb[53]  (.D(early_flags_lsb_Z[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[53]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_40 (.A(
        late_found_lsb_63_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[46]), .D(late_flags_lsb_Z[110]), .FCI(
        late_found_lsb_63_2_1_co0_19), .S(
        late_found_lsb_63_2_1_wmux_40_S), .Y(
        late_found_lsb_63_2_1_y5_2), .FCO(late_found_lsb_63_2_1_co1_19)
        );
    SLE \early_flags_lsb[113]  (.D(early_flags_lsb_Z[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[113]));
    CFG3 #( .INIT(8'h01) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_1_sqmuxa_1_0_a3_2  
        (.A(clkalign_curr_state_Z[1]), .B(N_533), .C(
        clkalign_curr_state_Z[0]), .Y(N_602_2));
    CFG4 #( .INIT(16'hECA0) )  
        \clkalign_curr_state_ns_5_0_.wait_cnt_3_o3[1]  (.A(N_659), .B(
        N_657), .C(clkalign_curr_state_Z[0]), .D(N_651), .Y(N_540));
    SLE \rst_cnt[4]  (.D(rst_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[4]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_28 (.A(
        early_found_msb_126_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[43]), .D(early_flags_msb_Z[107]), .FCI(
        early_found_msb_126_2_1_co0_13), .S(
        early_found_msb_126_2_1_wmux_28_S), .Y(
        early_found_msb_126_2_1_y5_1), .FCO(
        early_found_msb_126_2_1_co1_13));
    SLE \late_flags_lsb[21]  (.D(late_flags_lsb_Z[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[21]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[17])
        , .D(late_flags_msb_Z[81]), .FCI(late_found_msb_126_2_1_0_co1), 
        .S(late_found_msb_126_2_1_wmux_1_S), .Y(
        late_found_msb_126_2_1_y0_0), .FCO(
        late_found_msb_126_2_1_co0_0));
    SLE \late_flags_lsb[0]  (.D(late_flags_lsb_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_24 (.A(
        early_found_msb_63_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[34]), .D(early_flags_msb_Z[98]), .FCI(
        early_found_msb_63_2_1_co0_11), .S(
        early_found_msb_63_2_1_wmux_24_S), .Y(
        early_found_msb_63_2_1_y1_1), .FCO(
        early_found_msb_63_2_1_co1_11));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_21 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_126_2_1_co1_9), .S(
        early_found_lsb_126_2_1_wmux_21_S), .Y(
        early_found_lsb_126_2_1_wmux_21_Y), .FCO(
        early_found_lsb_126_2_1_co0_10));
    SLE \emflag_cnt[6]  (.D(emflag_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[19]), .D(early_flags_lsb_Z[83]), .FCI(
        early_found_lsb_126_2_1_co1_11), .S(
        early_found_lsb_126_2_1_wmux_25_S), .Y(
        early_found_lsb_126_2_1_y0_11), .FCO(
        early_found_lsb_126_2_1_co0_12));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_2 (.A(
        late_found_lsb_63_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[48]), .D(late_flags_lsb_Z[112]), .FCI(
        late_found_lsb_63_2_1_co0_0), .S(
        late_found_lsb_63_2_1_wmux_2_S), .Y(late_found_lsb_63_2_1_0_y3)
        , .FCO(late_found_lsb_63_2_1_co1_0));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_14 (.A(
        late_found_msb_126_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[53]), .D(late_flags_msb_Z[117]), .FCI(
        late_found_msb_126_2_1_co0_6), .S(
        late_found_msb_126_2_1_wmux_14_S), .Y(
        late_found_msb_126_2_1_y3_0), .FCO(
        late_found_msb_126_2_1_co1_6));
    SLE \early_late_start_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[5]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_14 (.A(
        early_found_msb_63_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[52]), .D(early_flags_msb_Z[116]), .FCI(
        early_found_msb_63_2_1_co0_6), .S(
        early_found_msb_63_2_1_wmux_14_S), .Y(
        early_found_msb_63_2_1_y3_0), .FCO(
        early_found_msb_63_2_1_co1_6));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[6])
        , .D(early_flags_lsb_Z[70]), .FCI(
        early_found_lsb_63_2_1_co1_16), .S(
        early_found_lsb_63_2_1_wmux_35_S), .Y(
        early_found_lsb_63_2_1_y0_15), .FCO(
        early_found_lsb_63_2_1_co0_17));
    SLE \early_flags_lsb[92]  (.D(early_flags_lsb_Z[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[92]));
    SLE \late_flags_msb[18]  (.D(late_flags_msb_Z[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[18]));
    ARI1 #( .INIT(20'h0CEC2) )  late_found_lsb_126_2_1_wmux_10 (.A(
        late_found_lsb_126_2_1_0_y21), .B(late_found_lsb_126_2_1_0_y9), 
        .C(emflag_cnt_Z[2]), .D(emflag_cnt_Z[1]), .FCI(
        late_found_lsb_126_2_1_co0_4), .S(
        late_found_lsb_126_2_1_wmux_10_S), .Y(
        late_found_lsb_126_2_1_y0_4), .FCO(
        late_found_lsb_126_2_1_co1_4));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_4 (.A(
        early_late_init_val_Z[4]), .B(early_late_nxt_val_Z[4]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_3_Z), .S(
        un2_sig_tapcnt_final_2_cry_4_S), .Y(
        un2_sig_tapcnt_final_2_cry_4_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_4_Z));
    SLE \rst_cnt[2]  (.D(rst_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[2]));
    SLE \late_flags_lsb[81]  (.D(late_flags_lsb_Z[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[81]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[2])
        , .D(early_flags_lsb_Z[66]), .FCI(
        early_found_lsb_63_2_1_co1_10), .S(
        early_found_lsb_63_2_1_wmux_23_S), .Y(
        early_found_lsb_63_2_1_y0_10), .FCO(
        early_found_lsb_63_2_1_co0_11));
    CFG2 #( .INIT(4'h2) )  \clkalign_curr_state_ns_5_0_.m35  (.A(N_30), 
        .B(N_127_mux), .Y(N_134_mux));
    SLE \late_flags_lsb[25]  (.D(late_flags_lsb_Z[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[25]));
    SLE calc_done (.D(calc_done_0_sqmuxa), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_17_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(calc_done_Z));
    CFG4 #( .INIT(16'hF088) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_1_sqmuxa_1_0_a3_RNIN2AC  
        (.A(N_643), .B(N_644), .C(tap_cnt_Z[7]), .D(
        clkalign_curr_state_1_sqmuxa_1), .Y(un1_early_flags_lsb14_i));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_16 (.A(
        late_found_msb_126_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[45]), .D(late_flags_msb_Z[109]), .FCI(
        late_found_msb_126_2_1_co0_7), .S(
        late_found_msb_126_2_1_wmux_16_S), .Y(
        late_found_msb_126_2_1_y5_0), .FCO(
        late_found_msb_126_2_1_co1_7));
    SLE \early_flags_lsb[127]  (.D(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[127]));
    SLE \early_flags_msb[127]  (.D(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[127]));
    SLE \late_flags_lsb[77]  (.D(late_flags_lsb_Z[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[77]));
    CFG4 #( .INIT(16'h0800) )  
        \clkalign_curr_state_ns_5_0_.clk_align_start6_0_a3  (.A(N_651), 
        .B(current_state_0), .C(clkalign_curr_state_Z[1]), .D(N_639), 
        .Y(clk_align_start6));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_7 
        (.A(early_late_end_val_Z[7]), .B(early_late_start_val_Z[7]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_6_Z), .S(
        early_late_start_end_val_status5_cry_7_S), .Y(
        early_late_start_end_val_status5_cry_7_Y), .FCO(
        early_late_start_end_val_status5));
    CFG2 #( .INIT(4'h4) )  
        \clkalign_curr_state_ns_5_0_.reset_dly_fg4_4  (.A(
        reset_dly_fg_Z), .B(rst_cnt_Z[8]), .Y(reset_dly_fg4_4));
    SLE \early_flags_msb[34]  (.D(early_flags_msb_Z[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[34]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_20 (.A(
        early_found_msb_126_2_1_y0_9), .B(early_found_msb_126_2_1_y3_0)
        , .C(early_found_msb_126_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_126_2_1_co0_9), .S(
        early_found_msb_126_2_1_wmux_20_S), .Y(
        early_found_msb_126_2_1_0_y21), .FCO(
        early_found_msb_126_2_1_co1_9));
    SLE \early_flags_lsb[60]  (.D(early_flags_lsb_Z[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[60]));
    SLE \sig_tapcnt_final_1[2]  (.D(sig_tapcnt_final_1_3_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[2]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_63_2_1_wmux_33 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_63_2_1_co1_15), .S(
        late_found_msb_63_2_1_wmux_33_S), .Y(
        late_found_msb_63_2_1_wmux_33_Y), .FCO(
        late_found_msb_63_2_1_co0_16));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_33 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_126_2_1_co1_15), .S(
        late_found_lsb_126_2_1_wmux_33_S), .Y(
        late_found_lsb_126_2_1_wmux_33_Y), .FCO(
        late_found_lsb_126_2_1_co0_16));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[23]), .D(early_flags_msb_Z[87]), .FCI(
        early_found_msb_126_2_1_co1_17), .S(
        early_found_msb_126_2_1_wmux_37_S), .Y(
        early_found_msb_126_2_1_y0_16), .FCO(
        early_found_msb_126_2_1_co0_18));
    SLE \early_flags_msb[82]  (.D(early_flags_msb_Z[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[82]));
    SLE \early_flags_lsb[75]  (.D(early_flags_lsb_Z[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[75]));
    SLE \late_flags_lsb[85]  (.D(late_flags_lsb_Z[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[85]));
    SLE early_or_late_found_msb_d (.D(early_or_late_found_msb_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_or_late_found_msb_d_Z));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_16 (.A(
        early_found_lsb_126_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[45]), .D(early_flags_lsb_Z[109]), .FCI(
        early_found_lsb_126_2_1_co0_7), .S(
        early_found_lsb_126_2_1_wmux_16_S), .Y(
        early_found_lsb_126_2_1_y5_0), .FCO(
        early_found_lsb_126_2_1_co1_7));
    CFG4 #( .INIT(16'h1302) )  \clkalign_curr_state_ns_5_0_.m117  (.A(
        clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[3]), .C(
        N_131_mux), .D(clkalign_curr_state_Z[4]), .Y(N_118));
    SLE \early_flags_lsb[32]  (.D(early_flags_lsb_Z[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[32]));
    SLE \early_late_init_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[6]));
    ARI1 #( .INIT(20'h555AA) )  un3_sig_tapcnt_final_1_cry_5 (.A(
        early_late_end_val_Z[5]), .B(early_late_start_val_Z[5]), .C(
        GND), .D(GND), .FCI(un3_sig_tapcnt_final_1_cry_4_Z), .S(
        un3_sig_tapcnt_final_1_cry_5_S), .Y(
        un3_sig_tapcnt_final_1_cry_5_Y), .FCO(
        un3_sig_tapcnt_final_1_cry_5_Z));
    SLE \late_flags_msb[61]  (.D(late_flags_msb_Z[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[61]));
    SLE \late_flags_lsb[1]  (.D(late_flags_lsb_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[1]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_126_2_1_wmux_19 (.A(
        early_found_lsb_126_2_1_y7_0), .B(early_found_lsb_126_2_1_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_126_2_1_co1_8), .S(
        early_found_lsb_126_2_1_wmux_19_S), .Y(
        early_found_lsb_126_2_1_y0_9), .FCO(
        early_found_lsb_126_2_1_co0_9));
    CFG4 #( .INIT(16'h0001) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_nxt_set14_3_i_a3_RNI3H371  
        (.A(N_637), .B(N_639), .C(N_549), .D(N_620), .Y(N_517_i));
    SLE \early_flags_msb[22]  (.D(early_flags_msb_Z[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[22]));
    SLE \early_flags_msb[31]  (.D(early_flags_msb_Z[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[31]));
    SLE \early_flags_msb[67]  (.D(early_flags_msb_Z[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[67]));
    SLE \late_flags_msb[5]  (.D(late_flags_msb_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[5]));
    SLE \early_flags_lsb[20]  (.D(early_flags_lsb_Z[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[20]));
    SLE \early_flags_lsb[107]  (.D(early_flags_lsb_Z[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[107]));
    SLE \early_flags_msb[107]  (.D(early_flags_msb_Z[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[107]));
    SLE \early_flags_msb[116]  (.D(early_flags_msb_Z[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[116]));
    CFG3 #( .INIT(8'hBF) )  \clkalign_curr_state_ns_5_0_.tap_cnt9_i  (
        .A(tap_cnt9_i_0), .B(N_2979), .C(N_125_mux), .Y(N_490));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[20]), .D(early_flags_lsb_Z[84]), .FCI(
        early_found_lsb_63_2_1_co1_5), .S(
        early_found_lsb_63_2_1_wmux_13_S), .Y(
        early_found_lsb_63_2_1_y0_6), .FCO(
        early_found_lsb_63_2_1_co0_6));
    SLE \late_flags_lsb[66]  (.D(late_flags_lsb_Z[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[66]));
    CFG4 #( .INIT(16'h0001) )  
        \clkalign_curr_state_ns_5_0_.rx_trng_done_3_0_0_958_a2  (.A(
        wait_cnt_Z[1]), .B(wait_cnt_Z[0]), .C(clkalign_curr_state_Z[2])
        , .D(wait_cnt_Z[2]), .Y(N_2967));
    CFG4 #( .INIT(16'hC682) )  \clkalign_curr_state_ns_5_0_.m104  (.A(
        clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[2]), .C(
        m104_1_2), .D(N_97), .Y(N_105));
    SLE \late_flags_msb[65]  (.D(late_flags_msb_Z[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[65]));
    SLE \late_flags_lsb[63]  (.D(late_flags_lsb_Z[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[63]));
    SLE \early_flags_msb[36]  (.D(early_flags_msb_Z[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[36]));
    CFG4 #( .INIT(16'h8000) )  emflag_cnt_done (.A(emflag_cnt_Z[1]), 
        .B(emflag_cnt_Z[2]), .C(emflag_cnt_done_5_Z), .D(
        emflag_cnt_Z[6]), .Y(emflag_cnt_done_Z));
    SLE early_late_init_set (.D(clkalign_curr_state_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(early_late_init_set_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_37 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[23])
        , .D(late_flags_msb_Z[87]), .FCI(late_found_msb_126_2_1_co1_17)
        , .S(late_found_msb_126_2_1_wmux_37_S), .Y(
        late_found_msb_126_2_1_y0_16), .FCO(
        late_found_msb_126_2_1_co0_18));
    SLE \late_flags_lsb[74]  (.D(late_flags_lsb_Z[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[74]));
    CFG4 #( .INIT(16'h5155) )  \clkalign_curr_state_ns_5_0_.m21  (.A(
        clkalign_curr_state_Z[4]), .B(N_19_i), .C(rx_err_Z), .D(
        calc_done_Z), .Y(N_139_mux));
    CFG4 #( .INIT(16'h7737) )  \clkalign_curr_state_ns_5_0_.m49  (.A(
        emflag_cnt_done_d_Z), .B(clkalign_curr_state_Z[0]), .C(
        no_early_and_late_found_Z), .D(early_or_late_found_Z), .Y(
        N_130_mux));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_5 (.A(
        early_late_init_val_Z[5]), .B(early_late_nxt_val_Z[5]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_4_Z), .S(
        un2_sig_tapcnt_final_2_cry_5_S), .Y(
        un2_sig_tapcnt_final_2_cry_5_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_5_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[7]  (.A(VCC), .B(
        rst_cnt_Z[7]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[6]), .S(
        rst_cnt_s[7]), .Y(rst_cnt_cry_Y[7]), .FCO(rst_cnt_cry_Z[7]));
    SLE \late_flags_msb[46]  (.D(late_flags_msb_Z[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[46]));
    SLE \late_flags_msb[43]  (.D(late_flags_msb_Z[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[43]));
    SLE \late_flags_msb[4]  (.D(late_flags_msb_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[4]));
    ARI1 #( .INIT(20'h0EA4A) )  late_found_lsb_126_2_1_wmux_9 (.A(
        late_found_lsb_126_2_1_0_y45), .B(late_found_lsb_126_2_1_y0_4), 
        .C(late_found_lsb_126_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        late_found_lsb_126_2_1_co1_3), .S(
        late_found_lsb_126_2_1_wmux_9_S), .Y(N_2094), .FCO(
        late_found_lsb_126_2_1_co0_4));
    SLE \late_flags_lsb[92]  (.D(late_flags_lsb_Z[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[92]));
    SLE no_early_and_late_found_lsb_d (.D(
        no_early_and_late_found_lsb_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(no_early_and_late_found_lsb_d_Z));
    SLE \late_flags_msb[119]  (.D(late_flags_msb_Z[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[119]));
    SLE \late_flags_msb[103]  (.D(late_flags_msb_Z[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[103]));
    CFG3 #( .INIT(8'h40) )  
        \clkalign_curr_state_ns_5_0_.start_trng_fg6  (.A(timeout_fg), 
        .B(current_state_0), .C(reset_dly_fg_Z), .Y(start_trng_fg6));
    CFG2 #( .INIT(4'h8) )  \clkalign_curr_state_ns_5_0_.m26  (.A(
        clkalign_curr_state81), .B(N_125_mux), .Y(N_27));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_18 (.A(
        late_found_msb_63_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[60]), .D(late_flags_msb_Z[124]), .FCI(
        late_found_msb_63_2_1_co0_8), .S(
        late_found_msb_63_2_1_wmux_18_S), .Y(
        late_found_msb_63_2_1_y7_0), .FCO(late_found_msb_63_2_1_co1_8));
    SLE \early_flags_msb[38]  (.D(early_flags_msb_Z[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[38]));
    SLE \late_flags_msb[19]  (.D(late_flags_msb_Z[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[19]));
    SLE \early_flags_lsb[95]  (.D(early_flags_lsb_Z[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[95]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_0 (.A(
        early_found_lsb_63_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[32]), .D(early_flags_lsb_Z[96]), .FCI(
        early_found_lsb_63_2_1_0_co0), .S(
        early_found_lsb_63_2_1_wmux_0_S), .Y(
        early_found_lsb_63_2_1_0_y1), .FCO(
        early_found_lsb_63_2_1_0_co1));
    CFG3 #( .INIT(8'hB8) )  \clkalign_curr_state_ns_5_0_.m82  (.A(N_30)
        , .B(clkalign_curr_state_Z[1]), .C(N_82_i), .Y(N_83));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_38 (.A(
        late_found_lsb_63_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[54]), .D(late_flags_lsb_Z[118]), .FCI(
        late_found_lsb_63_2_1_co0_18), .S(
        late_found_lsb_63_2_1_wmux_38_S), .Y(
        late_found_lsb_63_2_1_y3_2), .FCO(late_found_lsb_63_2_1_co1_18)
        );
    SLE \early_flags_msb[13]  (.D(early_flags_msb_Z[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[13]));
    SLE \late_flags_msb[36]  (.D(late_flags_msb_Z[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[36]));
    SLE \late_flags_msb[33]  (.D(late_flags_msb_Z[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[33]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_63_2_1_wmux_34 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_63_2_1_co0_16), .S(
        early_found_msb_63_2_1_wmux_34_S), .Y(
        early_found_msb_63_2_1_wmux_34_Y), .FCO(
        early_found_msb_63_2_1_co1_16));
    SLE \late_flags_msb[107]  (.D(late_flags_msb_Z[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[107]));
    SLE \early_flags_msb[50]  (.D(early_flags_msb_Z[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[50]));
    SLE \early_flags_msb[64]  (.D(early_flags_msb_Z[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[64]));
    SLE \late_flags_msb[86]  (.D(late_flags_msb_Z[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[86]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[1])
        , .D(early_flags_lsb_Z[65]), .FCI(VCC), .S(
        early_found_lsb_126_2_1_0_wmux_S), .Y(
        early_found_lsb_126_2_1_0_y0), .FCO(
        early_found_lsb_126_2_1_0_co0));
    CFG2 #( .INIT(4'hD) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final20_i_o3  (.A(
        early_late_init_and_nxt_set_Z), .B(tapcnt_final_2_status_Z), 
        .Y(N_552_i));
    SLE \late_flags_msb[83]  (.D(late_flags_msb_Z[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[83]));
    SLE \late_flags_msb[21]  (.D(late_flags_msb_Z[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[21]));
    SLE \early_flags_msb[85]  (.D(early_flags_msb_Z[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[85]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_6 (.A(
        early_found_lsb_63_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[56]), .D(early_flags_lsb_Z[120]), .FCI(
        early_found_lsb_63_2_1_co0_2), .S(
        early_found_lsb_63_2_1_wmux_6_S), .Y(
        early_found_lsb_63_2_1_0_y7), .FCO(
        early_found_lsb_63_2_1_co1_2));
    SLE \early_flags_msb[49]  (.D(early_flags_msb_Z[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[49]));
    CFG4 #( .INIT(16'h0001) )  sig_tapcnt_final_210_4 (.A(
        early_late_nxt_val_Z[7]), .B(early_late_nxt_val_Z[6]), .C(
        early_late_nxt_val_Z[4]), .D(early_late_nxt_val_Z[1]), .Y(
        sig_tapcnt_final_210_4_Z));
    SLE \clkalign_curr_state[5]  (.D(clkalign_curr_state_ns[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(clkalign_curr_state_Z[5]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_28 (.A(
        late_found_msb_63_2_1_y0_12), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[42]), .D(late_flags_msb_Z[106]), .FCI(
        late_found_msb_63_2_1_co0_13), .S(
        late_found_msb_63_2_1_wmux_28_S), .Y(
        late_found_msb_63_2_1_y5_1), .FCO(late_found_msb_63_2_1_co1_13)
        );
    SLE \early_flags_lsb[35]  (.D(early_flags_lsb_Z[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[35]));
    SLE \late_flags_msb[78]  (.D(late_flags_msb_Z[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[78]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[0]), 
        .D(late_flags_lsb_Z[64]), .FCI(VCC), .S(
        late_found_lsb_63_2_1_0_wmux_S), .Y(late_found_lsb_63_2_1_0_y0)
        , .FCO(late_found_lsb_63_2_1_0_co0));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_18 (.A(
        early_found_lsb_126_2_1_y0_8), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[61]), .D(early_flags_lsb_Z[125]), .FCI(
        early_found_lsb_126_2_1_co0_8), .S(
        early_found_lsb_126_2_1_wmux_18_S), .Y(
        early_found_lsb_126_2_1_y7_0), .FCO(
        early_found_lsb_126_2_1_co1_8));
    ARI1 #( .INIT(20'h4AA00) )  \timeout_cnt_s[7]  (.A(VCC), .B(
        timeout_cnt_Z[7]), .C(GND), .D(GND), .FCI(timeout_cnt_cry_Z[6])
        , .S(timeout_cnt_s_Z[7]), .Y(timeout_cnt_s_Y[7]), .FCO(
        timeout_cnt_s_FCO[7]));
    SLE \sig_tapcnt_final_2[5]  (.D(sig_tapcnt_final_2_3_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[5]));
    SLE \late_flags_lsb[125]  (.D(late_flags_lsb_Z[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[125]));
    SLE \early_flags_msb[25]  (.D(early_flags_msb_Z[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[25]));
    SLE \late_flags_lsb[101]  (.D(late_flags_lsb_Z[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[101]));
    SLE \early_flags_msb[61]  (.D(early_flags_msb_Z[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[61]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[15])
        , .D(late_flags_lsb_Z[79]), .FCI(late_found_lsb_126_2_1_co1_18)
        , .S(late_found_lsb_126_2_1_wmux_39_S), .Y(
        late_found_lsb_126_2_1_y0_17), .FCO(
        late_found_lsb_126_2_1_co0_19));
    SLE \late_flags_msb[25]  (.D(late_flags_msb_Z[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[25]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[5]  (.A(VCC), .B(
        rst_cnt_Z[5]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[4]), .S(
        rst_cnt_s[5]), .Y(rst_cnt_cry_Y[5]), .FCO(rst_cnt_cry_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[8])
        , .D(early_flags_lsb_Z[72]), .FCI(early_found_lsb_63_2_1_co1_0)
        , .S(early_found_lsb_63_2_1_wmux_3_S), .Y(
        early_found_lsb_63_2_1_y0_1), .FCO(
        early_found_lsb_63_2_1_co0_1));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_s[9]  (.A(VCC), .B(
        rst_cnt_Z[9]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[8]), .S(
        rst_cnt_s_Z[9]), .Y(rst_cnt_s_Y[9]), .FCO(rst_cnt_s_FCO[9]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_42 (.A(
        early_found_msb_126_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[63]), .D(early_flags_msb_Z[127]), .FCI(
        early_found_msb_126_2_1_co0_20), .S(
        early_found_msb_126_2_1_wmux_42_S), .Y(
        early_found_msb_126_2_1_y7_2), .FCO(
        early_found_msb_126_2_1_co1_20));
    SLE \early_flags_msb[66]  (.D(early_flags_msb_Z[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[66]));
    CFG4 #( .INIT(16'hEDFF) )  
        \clkalign_curr_state_ns_5_0_.tap_cnt9_i_0  (.A(
        clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[5]), .C(
        clkalign_curr_state_Z[1]), .D(clkalign_curr_state_Z[0]), .Y(
        tap_cnt9_i_0));
    SLE \early_flags_lsb[43]  (.D(early_flags_lsb_Z[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[43]));
    SLE early_not_found_lsb_d (.D(early_found_lsb_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_not_found_lsb_d_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_25 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[18]), .D(early_flags_msb_Z[82]), .FCI(
        early_found_msb_63_2_1_co1_11), .S(
        early_found_msb_63_2_1_wmux_25_S), .Y(
        early_found_msb_63_2_1_y0_11), .FCO(
        early_found_msb_63_2_1_co0_12));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[1]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_2_S), 
        .Y(sig_tapcnt_final_1_3_Z[1]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[25]), .D(early_flags_lsb_Z[89]), .FCI(
        early_found_lsb_126_2_1_co1_1), .S(
        early_found_lsb_126_2_1_wmux_5_S), .Y(
        early_found_lsb_126_2_1_y0_2), .FCO(
        early_found_lsb_126_2_1_co0_2));
    CFG3 #( .INIT(8'h27) )  late_found_msb_127_i (.A(emflag_cnt_Z[0]), 
        .B(N_2348), .C(N_2285), .Y(late_found_msb_i));
    CFG4 #( .INIT(16'hECCC) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_8_0_0  
        (.A(N_602_2), .B(N_622), .C(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), .D(N_2979), .Y(
        un1_clkalign_curr_state_0_sqmuxa_8_0_0));
    CFG4 #( .INIT(16'hFFFE) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_17_0  (.A(
        N_593), .B(clkalign_curr_state_d[27]), .C(N_585_i), .D(N_594), 
        .Y(un1_clkalign_curr_state_17_0));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_63_2_1_wmux_31 (.A(
        late_found_msb_63_2_1_y7_1), .B(late_found_msb_63_2_1_y5_1), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co1_14), .S(
        late_found_msb_63_2_1_wmux_31_S), .Y(
        late_found_msb_63_2_1_y0_14), .FCO(
        late_found_msb_63_2_1_co0_15));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[16])
        , .D(late_flags_msb_Z[80]), .FCI(late_found_msb_63_2_1_0_co1), 
        .S(late_found_msb_63_2_1_wmux_1_S), .Y(
        late_found_msb_63_2_1_y0_0), .FCO(late_found_msb_63_2_1_co0_0));
    SLE \late_flags_lsb[2]  (.D(late_flags_lsb_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[2]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[12]), .D(early_flags_msb_Z[76]), .FCI(
        early_found_msb_63_2_1_co1_6), .S(
        early_found_msb_63_2_1_wmux_15_S), .Y(
        early_found_msb_63_2_1_y0_7), .FCO(
        early_found_msb_63_2_1_co0_7));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[17]), .D(early_flags_lsb_Z[81]), .FCI(
        early_found_lsb_126_2_1_0_co1), .S(
        early_found_lsb_126_2_1_wmux_1_S), .Y(
        early_found_lsb_126_2_1_y0_0), .FCO(
        early_found_lsb_126_2_1_co0_0));
    SLE \late_flags_msb[96]  (.D(late_flags_msb_Z[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[96]));
    SLE \early_flags_msb[99]  (.D(early_flags_msb_Z[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[99]));
    SLE \late_flags_msb[93]  (.D(late_flags_msb_Z[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[93]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[8]), 
        .D(late_flags_lsb_Z[72]), .FCI(late_found_lsb_63_2_1_co1_0), 
        .S(late_found_lsb_63_2_1_wmux_3_S), .Y(
        late_found_lsb_63_2_1_y0_1), .FCO(late_found_lsb_63_2_1_co0_1));
    GND GND_Z (.Y(GND));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[2]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_3_S), 
        .Y(sig_tapcnt_final_2_3_Z[2]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[5])
        , .D(early_flags_msb_Z[69]), .FCI(
        early_found_msb_126_2_1_co1_4), .S(
        early_found_msb_126_2_1_wmux_11_S), .Y(
        early_found_msb_126_2_1_y0_5), .FCO(
        early_found_msb_126_2_1_co0_5));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[31])
        , .D(late_flags_msb_Z[95]), .FCI(late_found_msb_126_2_1_co1_19)
        , .S(late_found_msb_126_2_1_wmux_41_S), .Y(
        late_found_msb_126_2_1_y0_18), .FCO(
        late_found_msb_126_2_1_co0_20));
    CFG2 #( .INIT(4'h8) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_s5_0_a2_0  (
        .A(clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[0]), .Y(
        N_644));
    SLE \early_flags_msb[68]  (.D(early_flags_msb_Z[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[68]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_63_2_1_wmux_42 (.A(
        early_found_lsb_63_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[62]), .D(early_flags_lsb_Z[126]), .FCI(
        early_found_lsb_63_2_1_co0_20), .S(
        early_found_lsb_63_2_1_wmux_42_S), .Y(
        early_found_lsb_63_2_1_y7_2), .FCO(
        early_found_lsb_63_2_1_co1_20));
    SLE \early_flags_lsb[2]  (.D(early_flags_lsb_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[2]));
    CFG1 #( .INIT(2'h1) )  \rst_cnt_RNO[0]  (.A(rst_cnt_Z[0]), .Y(
        rst_cnt_s[0]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_6 (.A(
        late_found_lsb_126_2_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[57]), .D(late_flags_lsb_Z[121]), .FCI(
        late_found_lsb_126_2_1_co0_2), .S(
        late_found_lsb_126_2_1_wmux_6_S), .Y(
        late_found_lsb_126_2_1_0_y7), .FCO(
        late_found_lsb_126_2_1_co1_2));
    SLE \late_flags_lsb[97]  (.D(late_flags_lsb_Z[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[97]));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[0]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[0]), .D(GND), .FCI(
        tap_cnt_cry_cy), .S(tap_cnt_s[0]), .Y(tap_cnt_cry_Y[0]), .FCO(
        tap_cnt_cry_Z[0]));
    SLE \late_flags_lsb[16]  (.D(late_flags_lsb_Z[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[16]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_2 (.A(
        late_found_msb_63_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[48]), .D(late_flags_msb_Z[112]), .FCI(
        late_found_msb_63_2_1_co0_0), .S(
        late_found_msb_63_2_1_wmux_2_S), .Y(late_found_msb_63_2_1_0_y3)
        , .FCO(late_found_msb_63_2_1_co1_0));
    SLE \late_flags_lsb[13]  (.D(late_flags_lsb_Z[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[13]));
    SLE \late_flags_lsb[115]  (.D(late_flags_lsb_Z[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[115]));
    ARI1 #( .INIT(20'h0FA44) )  
        \clkalign_curr_state_ns_5_0_.m70_1_0_wmux  (.A(
        clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[3]), .C(
        N_46), .D(N_58), .FCI(VCC), .S(m70_1_0_wmux_S), .Y(m70_1_0_y0), 
        .FCO(m70_1_0_co0));
    CFG2 #( .INIT(4'h8) )  \clkalign_curr_state_ns_5_0_.m18  (.A(
        clkalign_curr_state_Z[0]), .B(N_125_mux), .Y(N_19_i));
    SLE \early_flags_msb[121]  (.D(early_flags_msb_Z[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[121]));
    CFG3 #( .INIT(8'h40) )  \clkalign_curr_state_ns_5_0_.m41  (.A(
        clkalign_curr_state_Z[4]), .B(start_trng_fg_Z), .C(
        clkalign_curr_state_Z[0]), .Y(N_128_mux));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.un1_internal_rst_en_2_0  (.A(
        clk_align_start6), .B(N_585_i), .Y(un1_internal_rst_en_2_0));
    SLE \sig_tapcnt_final_2[0]  (.D(sig_tapcnt_final_2_3_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[0]));
    CFG4 #( .INIT(16'hEE30) )  \clkalign_curr_state_ns_5_0_.m114_2  (
        .A(N_109), .B(clkalign_curr_state_Z[1]), .C(N_139_mux), .D(
        m114_2_1), .Y(N_115));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_21 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_126_2_1_co1_9), .S(
        late_found_msb_126_2_1_wmux_21_S), .Y(
        late_found_msb_126_2_1_wmux_21_Y), .FCO(
        late_found_msb_126_2_1_co0_10));
    SLE tapcnt_final_1_status (.D(sig_tapcnt_final_111_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_final_1_status_Z));
    SLE \late_flags_msb[79]  (.D(late_flags_msb_Z[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[79]));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_0 (.A(
        early_late_init_val_Z[0]), .B(early_late_nxt_val_Z[0]), .C(GND)
        , .D(GND), .FCI(GND), .S(un2_sig_tapcnt_final_2_cry_0_S), .Y(
        un2_sig_tapcnt_final_2_cry_0_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_0_Z));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_4 (.A(
        late_found_lsb_63_2_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[40]), .D(late_flags_lsb_Z[104]), .FCI(
        late_found_lsb_63_2_1_co0_1), .S(
        late_found_lsb_63_2_1_wmux_4_S), .Y(late_found_lsb_63_2_1_0_y5)
        , .FCO(late_found_lsb_63_2_1_co1_1));
    ARI1 #( .INIT(20'h0EA4A) )  early_found_msb_126_2_1_wmux_9 (.A(
        early_found_msb_126_2_1_0_y45), .B(
        early_found_msb_126_2_1_y0_4), .C(
        early_found_msb_126_2_1_0_y33), .D(emflag_cnt_Z[1]), .FCI(
        early_found_msb_126_2_1_co1_3), .S(
        early_found_msb_126_2_1_wmux_9_S), .Y(N_2221), .FCO(
        early_found_msb_126_2_1_co0_4));
    SLE early_late_init_nxt_val_status (.D(
        early_late_init_nxt_val_status5), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_late_init_nxt_val_status_Z));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_21 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_63_2_1_co1_9), .S(
        early_found_lsb_63_2_1_wmux_21_S), .Y(
        early_found_lsb_63_2_1_wmux_21_Y), .FCO(
        early_found_lsb_63_2_1_co0_10));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[3]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_4_S), 
        .Y(sig_tapcnt_final_2_3_Z[3]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_22 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_msb_126_2_1_co0_10), .S(
        early_found_msb_126_2_1_wmux_22_S), .Y(
        early_found_msb_126_2_1_wmux_22_Y), .FCO(
        early_found_msb_126_2_1_co1_10));
    SLE \late_flags_lsb[71]  (.D(late_flags_lsb_Z[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[71]));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_42 (.A(
        early_found_lsb_126_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[63]), .D(early_flags_lsb_Z[127]), .FCI(
        early_found_lsb_126_2_1_co0_20), .S(
        early_found_lsb_126_2_1_wmux_42_S), .Y(
        early_found_lsb_126_2_1_y7_2), .FCO(
        early_found_lsb_126_2_1_co1_20));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[24]), .D(early_flags_lsb_Z[88]), .FCI(
        early_found_lsb_63_2_1_co1_1), .S(
        early_found_lsb_63_2_1_wmux_5_S), .Y(
        early_found_lsb_63_2_1_y0_2), .FCO(
        early_found_lsb_63_2_1_co0_2));
    SLE \early_flags_msb[32]  (.D(early_flags_msb_Z[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[32]));
    SLE \early_flags_msb[101]  (.D(early_flags_msb_Z[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[101]));
    CFG4 #( .INIT(16'h8000) )  
        \clkalign_curr_state_ns_5_0_.reset_dly_fg4_8  (.A(rst_cnt_Z[9])
        , .B(rst_cnt_Z[7]), .C(rst_cnt_Z[6]), .D(reset_dly_fg4_6), .Y(
        reset_dly_fg4_8));
    SLE \late_flags_lsb[94]  (.D(late_flags_lsb_Z[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[94]));
    SLE early_late_nxt_set (.D(clkalign_curr_state_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(N_517_i), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_late_nxt_set_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[9]), 
        .D(late_flags_msb_Z[73]), .FCI(late_found_msb_126_2_1_co1_0), 
        .S(late_found_msb_126_2_1_wmux_3_S), .Y(
        late_found_msb_126_2_1_y0_1), .FCO(
        late_found_msb_126_2_1_co0_1));
    CFG3 #( .INIT(8'h27) )  early_found_lsb_127_i (.A(emflag_cnt_Z[0]), 
        .B(N_1967), .C(N_1904), .Y(early_found_lsb_i));
    SLE \early_flags_msb[4]  (.D(early_flags_msb_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[4]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[20])
        , .D(late_flags_lsb_Z[84]), .FCI(late_found_lsb_63_2_1_co1_5), 
        .S(late_found_lsb_63_2_1_wmux_13_S), .Y(
        late_found_lsb_63_2_1_y0_6), .FCO(late_found_lsb_63_2_1_co0_6));
    SLE \late_flags_lsb[60]  (.D(late_flags_lsb_Z[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[60]));
    SLE rx_trng_done (.D(N_2967), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(un1_clkalign_curr_state_1_0), .ALn(current_state_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_trng_done_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_39 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[15]), .D(early_flags_msb_Z[79]), .FCI(
        early_found_msb_126_2_1_co1_18), .S(
        early_found_msb_126_2_1_wmux_39_S), .Y(
        early_found_msb_126_2_1_y0_17), .FCO(
        early_found_msb_126_2_1_co0_19));
    CFG4 #( .INIT(16'h5557) )  \clkalign_curr_state_ns_5_0_.m91  (.A(
        clkalign_curr_state_Z[4]), .B(current_state_0), .C(
        clkalign_curr_state_Z[0]), .D(clkalign_curr_state_Z[1]), .Y(
        N_131_mux));
    SLE \early_flags_msb[115]  (.D(early_flags_msb_Z[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[115]));
    CFG4 #( .INIT(16'h3313) )  \clkalign_curr_state_ns_5_0_.m80  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), .C(
        N_78), .D(clkalign_curr_state_Z[4]), .Y(N_143_mux));
    SLE \late_flags_lsb[75]  (.D(late_flags_lsb_Z[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[75]));
    SLE \early_flags_lsb[108]  (.D(early_flags_lsb_Z[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[108]));
    CFG4 #( .INIT(16'hFFEA) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_8_0  
        (.A(N_643), .B(N_526), .C(N_642), .D(
        un1_clkalign_curr_state_0_sqmuxa_8_0_0), .Y(
        un1_clkalign_curr_state_0_sqmuxa_8_0));
    SLE \late_flags_lsb[3]  (.D(late_flags_lsb_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[3]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_34 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_msb_126_2_1_co0_16), .S(
        late_found_msb_126_2_1_wmux_34_S), .Y(
        late_found_msb_126_2_1_wmux_34_Y), .FCO(
        late_found_msb_126_2_1_co1_16));
    SLE \late_flags_lsb[107]  (.D(late_flags_lsb_Z[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[107]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_30 (.A(
        late_found_lsb_126_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[59]), .D(late_flags_lsb_Z[123]), .FCI(
        late_found_lsb_126_2_1_co0_14), .S(
        late_found_lsb_126_2_1_wmux_30_S), .Y(
        late_found_lsb_126_2_1_y7_1), .FCO(
        late_found_lsb_126_2_1_co1_14));
    SLE \late_flags_msb[40]  (.D(late_flags_msb_Z[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[40]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_63_2_1_wmux_43 (.A(
        late_found_msb_63_2_1_y7_2), .B(late_found_msb_63_2_1_y5_2), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_63_2_1_co1_20), .S(
        late_found_msb_63_2_1_wmux_43_S), .Y(
        late_found_msb_63_2_1_y0_19), .FCO(
        late_found_msb_63_2_1_co0_21));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[6])
        , .D(early_flags_msb_Z[70]), .FCI(
        early_found_msb_63_2_1_co1_16), .S(
        early_found_msb_63_2_1_wmux_35_S), .Y(
        early_found_msb_63_2_1_y0_15), .FCO(
        early_found_msb_63_2_1_co0_17));
    SLE \emflag_cnt[3]  (.D(emflag_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[3]));
    SLE early_late_start_and_end_set (.D(
        early_late_start_and_end_set5_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_late_start_and_end_set_Z));
    SLE \early_flags_lsb[67]  (.D(early_flags_lsb_Z[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[67]));
    CFG3 #( .INIT(8'hD7) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_end_set12_3_i_0  (
        .A(clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[4]), .C(
        clkalign_curr_state_Z[3]), .Y(un1_early_late_end_set12_3_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[1]  (.A(VCC), .B(
        rst_cnt_Z[1]), .C(GND), .D(GND), .FCI(rst_cnt_s_1133_FCO), .S(
        rst_cnt_s[1]), .Y(rst_cnt_cry_Y[1]), .FCO(rst_cnt_cry_Z[1]));
    SLE \early_flags_lsb[89]  (.D(early_flags_lsb_Z[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[89]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_36 (.A(
        late_found_msb_126_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[39]), .D(late_flags_msb_Z[103]), .FCI(
        late_found_msb_126_2_1_co0_17), .S(
        late_found_msb_126_2_1_wmux_36_S), .Y(
        late_found_msb_126_2_1_y1_2), .FCO(
        late_found_msb_126_2_1_co1_17));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_34 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_126_2_1_co0_16), .S(
        early_found_lsb_126_2_1_wmux_34_S), .Y(
        early_found_lsb_126_2_1_wmux_34_Y), .FCO(
        early_found_lsb_126_2_1_co1_16));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[4])
        , .D(early_flags_lsb_Z[68]), .FCI(early_found_lsb_63_2_1_co1_4)
        , .S(early_found_lsb_63_2_1_wmux_11_S), .Y(
        early_found_lsb_63_2_1_y0_5), .FCO(
        early_found_lsb_63_2_1_co0_5));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[1]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[1]), .D(early_late_init_val_Z[1]), .Y(
        tapcnt_final_11_iv_1[1]));
    CFG4 #( .INIT(16'h40FB) )  \clkalign_curr_state_ns_5_0_.m96  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[4]), .C(
        N_61), .D(m96_1_0), .Y(N_97));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_63_2_1_wmux_0 (.A(
        late_found_lsb_63_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[32]), .D(late_flags_lsb_Z[96]), .FCI(
        late_found_lsb_63_2_1_0_co0), .S(
        late_found_lsb_63_2_1_wmux_0_S), .Y(late_found_lsb_63_2_1_0_y1)
        , .FCO(late_found_lsb_63_2_1_0_co1));
    SLE \early_flags_lsb[111]  (.D(early_flags_lsb_Z[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[111]));
    SLE \early_flags_msb[73]  (.D(early_flags_msb_Z[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[73]));
    SLE \emflag_cnt[2]  (.D(emflag_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(emflag_cnt_Z[2]));
    CFG3 #( .INIT(8'h35) )  \clkalign_curr_state_ns_5_0_.m54_1_2  (.A(
        tapcnt_final_2_status_Z), .B(tapcnt_final_1_status_Z), .C(
        early_late_start_and_end_set_Z), .Y(m54_1_2));
    CFG4 #( .INIT(16'hFFAB) )  
        \clkalign_curr_state_ns_5_0_.emflag_cnt10_i_3_RNIEGLP  (.A(
        clkalign_curr_state_s9_0_a3), .B(emflag_cnt10_i_3), .C(
        emflag_cnt_done_d_Z), .D(timeout_cnte), .Y(emflag_cnte));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_126_2_1_wmux_7 (.A(
        early_found_lsb_126_2_1_0_y7), .B(early_found_lsb_126_2_1_0_y5)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_126_2_1_co1_2), .S(
        early_found_lsb_126_2_1_wmux_7_S), .Y(
        early_found_lsb_126_2_1_y0_3), .FCO(
        early_found_lsb_126_2_1_co0_3));
    CFG4 #( .INIT(16'h0004) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_nxt_set14_3_i_a3  
        (.A(emflag_cnt_done_d_Z), .B(clkalign_curr_state_Z[4]), .C(
        early_or_late_found_Z), .D(no_early_and_late_found_Z), .Y(
        N_620));
    CFG3 #( .INIT(8'h48) )  \clkalign_curr_state_ns_5_0_.N_2935_i  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), .C(
        clkalign_curr_state_Z[0]), .Y(N_2935_i));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_126_2_1_wmux_43 (.A(
        late_found_msb_126_2_1_y7_2), .B(late_found_msb_126_2_1_y5_2), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co1_20), .S(
        late_found_msb_126_2_1_wmux_43_S), .Y(
        late_found_msb_126_2_1_y0_19), .FCO(
        late_found_msb_126_2_1_co0_21));
    SLE \late_flags_msb[30]  (.D(late_flags_msb_Z[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[30]));
    SLE \early_flags_lsb[122]  (.D(early_flags_lsb_Z[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[122]));
    SLE \late_flags_msb[3]  (.D(late_flags_msb_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[3]));
    SLE \late_flags_msb[1]  (.D(late_flags_msb_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[1]));
    SLE \early_flags_lsb[27]  (.D(early_flags_lsb_Z[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[27]));
    CFG2 #( .INIT(4'h2) )  \clkalign_curr_state_ns_5_0_.m3  (.A(
        clkalign_curr_state_Z[0]), .B(N_125_mux), .Y(N_4));
    CFG3 #( .INIT(8'hFE) )  
        \clkalign_curr_state_ns_5_0_.emflag_cnt10_i_3  (.A(
        emflag_cnt10_i_1), .B(N_657), .C(emflag_cnt10_i_0), .Y(
        emflag_cnt10_i_3));
    SLE \late_flags_lsb[46]  (.D(late_flags_lsb_Z[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[46]));
    SLE \early_flags_msb[110]  (.D(early_flags_msb_Z[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[110]));
    SLE \late_flags_lsb[43]  (.D(late_flags_lsb_Z[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[43]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_2 (.A(
        early_found_msb_63_2_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[48]), .D(early_flags_msb_Z[112]), .FCI(
        early_found_msb_63_2_1_co0_0), .S(
        early_found_msb_63_2_1_wmux_2_S), .Y(
        early_found_msb_63_2_1_0_y3), .FCO(
        early_found_msb_63_2_1_co1_0));
    SLE \early_flags_msb[40]  (.D(early_flags_msb_Z[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[40]));
    CFG3 #( .INIT(8'hD8) )  late_found_lsb_127 (.A(emflag_cnt_Z[0]), 
        .B(N_2094), .C(N_2031), .Y(late_found_lsb));
    SLE \late_flags_msb[80]  (.D(late_flags_msb_Z[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[80]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_126_2_1_wmux_43 (.A(
        early_found_msb_126_2_1_y7_2), .B(early_found_msb_126_2_1_y5_2)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_126_2_1_co1_20), .S(
        early_found_msb_126_2_1_wmux_43_S), .Y(
        early_found_msb_126_2_1_y0_19), .FCO(
        early_found_msb_126_2_1_co0_21));
    SLE \wait_cnt[1]  (.D(wait_cnt_3[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(wait_cnt_Z[1]));
    SLE RX_CLK_ALIGN_DONE (.D(RX_CLK_ALIGN_DONE5), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE));
    SLE \early_late_nxt_val[7]  (.D(emflag_cnt_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[7]));
    CFG3 #( .INIT(8'hD8) )  early_found_lsb_127 (.A(emflag_cnt_Z[0]), 
        .B(N_1967), .C(N_1904), .Y(early_found_lsb));
    SLE \early_flags_msb[109]  (.D(early_flags_msb_Z[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[109]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[16]), .D(early_flags_msb_Z[80]), .FCI(
        early_found_msb_63_2_1_0_co1), .S(
        early_found_msb_63_2_1_wmux_1_S), .Y(
        early_found_msb_63_2_1_y0_0), .FCO(
        early_found_msb_63_2_1_co0_0));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_0 (.A(
        late_found_msb_63_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[32]), .D(late_flags_msb_Z[96]), .FCI(
        late_found_msb_63_2_1_0_co0), .S(
        late_found_msb_63_2_1_wmux_0_S), .Y(late_found_msb_63_2_1_0_y1)
        , .FCO(late_found_msb_63_2_1_0_co1));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_22 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_126_2_1_co0_10), .S(
        early_found_lsb_126_2_1_wmux_22_S), .Y(
        early_found_lsb_126_2_1_wmux_22_Y), .FCO(
        early_found_lsb_126_2_1_co1_10));
    SLE \late_flags_lsb[52]  (.D(late_flags_lsb_Z[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[52]));
    SLE \early_flags_lsb[102]  (.D(early_flags_lsb_Z[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[102]));
    CFG2 #( .INIT(4'hD) )  \clkalign_curr_state_ns_5_0_.N_2924_i  (.A(
        N_125_mux), .B(clkalign_curr_state_Z[3]), .Y(N_2924_i));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[3]), 
        .D(late_flags_msb_Z[67]), .FCI(late_found_msb_126_2_1_co1_10), 
        .S(late_found_msb_126_2_1_wmux_23_S), .Y(
        late_found_msb_126_2_1_y0_10), .FCO(
        late_found_msb_126_2_1_co0_11));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[5]), 
        .D(late_flags_msb_Z[69]), .FCI(late_found_msb_126_2_1_co1_4), 
        .S(late_found_msb_126_2_1_wmux_11_S), .Y(
        late_found_msb_126_2_1_y0_5), .FCO(
        late_found_msb_126_2_1_co0_5));
    SLE \late_flags_msb[120]  (.D(late_flags_msb_Z[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[120]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[27])
        , .D(late_flags_msb_Z[91]), .FCI(late_found_msb_126_2_1_co1_13)
        , .S(late_found_msb_126_2_1_wmux_29_S), .Y(
        late_found_msb_126_2_1_y0_13), .FCO(
        late_found_msb_126_2_1_co0_14));
    CFG4 #( .INIT(16'h0602) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_nxt_set14_1_0  (.A(
        clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[4]), .C(
        N_549), .D(N_653), .Y(un1_early_late_nxt_set14_1_0));
    SLE \early_flags_msb[62]  (.D(early_flags_msb_Z[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[62]));
    SLE \early_flags_msb[35]  (.D(early_flags_msb_Z[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[35]));
    SLE reset_dly_fg (.D(VCC), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(reset_dly_fg4), .ALn(current_state_0), .ADn(VCC), .SLn(VCC)
        , .SD(GND), .LAT(GND), .Q(reset_dly_fg_Z));
    SLE \early_late_nxt_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_nxt_set14_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_nxt_val_Z[1]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_lsb_126_2_1_wmux_7 (.A(
        late_found_lsb_126_2_1_0_y7), .B(late_found_lsb_126_2_1_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co1_2), .S(
        late_found_lsb_126_2_1_wmux_7_S), .Y(
        late_found_lsb_126_2_1_y0_3), .FCO(
        late_found_lsb_126_2_1_co0_3));
    SLE \early_flags_lsb[64]  (.D(early_flags_lsb_Z[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[64]));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_2_3[1]  (.A(
        sig_tapcnt_final_210_Z), .B(un2_sig_tapcnt_final_2_cry_2_S), 
        .Y(sig_tapcnt_final_2_3_Z[1]));
    SLE \late_flags_lsb[36]  (.D(late_flags_lsb_Z[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[36]));
    SLE \sig_tapcnt_final_1[4]  (.D(sig_tapcnt_final_1_3_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[4]));
    CFG2 #( .INIT(4'h2) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_0_sqmuxa_4_0_a2  
        (.A(N_125_mux), .B(clkalign_curr_state_Z[2]), .Y(N_642));
    SLE \late_flags_lsb[33]  (.D(late_flags_lsb_Z[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[33]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_63_2_1_wmux_42 (.A(
        early_found_msb_63_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[62]), .D(early_flags_msb_Z[126]), .FCI(
        early_found_msb_63_2_1_co0_20), .S(
        early_found_msb_63_2_1_wmux_42_S), .Y(
        early_found_msb_63_2_1_y7_2), .FCO(
        early_found_msb_63_2_1_co1_20));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_0[1]  (.A(
        early_late_start_end_val_status_Z), .B(tapcnt_final_0_sqmuxa_1)
        , .C(sig_tapcnt_final_1_Z[1]), .D(early_late_start_val_Z[1]), 
        .Y(tapcnt_final_11_iv_0[1]));
    SLE \early_flags_lsb[109]  (.D(early_flags_lsb_Z[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[109]));
    SLE \early_late_end_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[3]));
    CFG2 #( .INIT(4'h4) )  \sig_tapcnt_final_1_3[4]  (.A(
        sig_tapcnt_final_111_Z), .B(un3_sig_tapcnt_final_1_cry_5_S), 
        .Y(sig_tapcnt_final_1_3_Z[4]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[0]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[0]), .D(early_late_init_val_Z[0]), .Y(
        tapcnt_final_11_iv_1[0]));
    SLE \late_flags_msb[121]  (.D(late_flags_msb_Z[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[121]));
    SLE RX_CLK_ALIGN_DONE_rep (.D(RX_CLK_ALIGN_DONE5), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(RX_CLK_ALIGN_DONE_rep_Z));
    SLE \sig_tapcnt_final_1[5]  (.D(sig_tapcnt_final_1_3_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_1_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[29]), .D(early_flags_msb_Z[93]), .FCI(
        early_found_msb_126_2_1_co1_7), .S(
        early_found_msb_126_2_1_wmux_17_S), .Y(
        early_found_msb_126_2_1_y0_8), .FCO(
        early_found_msb_126_2_1_co0_8));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[1]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[1]), .D(GND), .FCI(
        emflag_cnt_cry_Z[0]), .S(emflag_cnt_s[1]), .Y(
        emflag_cnt_cry_Y[1]), .FCO(emflag_cnt_cry_Z[1]));
    SLE \early_flags_msb[90]  (.D(early_flags_msb_Z[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[90]));
    SLE \early_flags_msb[57]  (.D(early_flags_msb_Z[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[57]));
    SLE \early_flags_lsb[61]  (.D(early_flags_lsb_Z[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[61]));
    SLE \tapcnt_final[6]  (.D(tapcnt_final_11[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[6]));
    SLE \early_flags_lsb[24]  (.D(early_flags_lsb_Z[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[24]));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNIL33I5[6]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[6]), 
        .D(GND), .FCI(tapcnt_offset_cry[5]), .S(tapcnt_offset_s[6]), 
        .Y(tapcnt_offset_RNIL33I5_Y[6]), .FCO(tapcnt_offset_cry[6]));
    CFG4 #( .INIT(16'hCCCA) )  \clkalign_curr_state_ns_5_0_.m54  (.A(
        emflag_cnt_done_d_Z), .B(m54_1_2), .C(
        early_late_init_and_nxt_set_Z), .D(
        early_late_start_and_end_set_Z), .Y(N_55));
    SLE \late_flags_msb[90]  (.D(late_flags_msb_Z[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[90]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_44 (.A(
        late_found_lsb_126_2_1_y0_19), .B(late_found_lsb_126_2_1_y3_2), 
        .C(late_found_lsb_126_2_1_y1_2), .D(emflag_cnt_Z[3]), .FCI(
        late_found_lsb_126_2_1_co0_21), .S(
        late_found_lsb_126_2_1_wmux_44_S), .Y(
        late_found_lsb_126_2_1_0_y45), .FCO(
        late_found_lsb_126_2_1_co1_21));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[9])
        , .D(early_flags_msb_Z[73]), .FCI(
        early_found_msb_126_2_1_co1_0), .S(
        early_found_msb_126_2_1_wmux_3_S), .Y(
        early_found_msb_126_2_1_y0_1), .FCO(
        early_found_msb_126_2_1_co0_1));
    SLE \early_flags_lsb[124]  (.D(early_flags_lsb_Z[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[124]));
    SLE \tapcnt_final[1]  (.D(tapcnt_final_11[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[1]));
    SLE \early_flags_lsb[66]  (.D(early_flags_lsb_Z[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[66]));
    SLE \cnt[1]  (.D(N_554_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(VCC), .ALn(current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND)
        , .LAT(GND), .Q(cnt_Z[1]));
    SLE early_not_found_msb_d (.D(early_found_msb_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_not_found_msb_d_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[1]), 
        .D(late_flags_msb_Z[65]), .FCI(VCC), .S(
        late_found_msb_126_2_1_0_wmux_S), .Y(
        late_found_msb_126_2_1_0_y0), .FCO(
        late_found_msb_126_2_1_0_co0));
    SLE \early_flags_lsb[21]  (.D(early_flags_lsb_Z[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[21]));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_126_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[3])
        , .D(early_flags_msb_Z[67]), .FCI(
        early_found_msb_126_2_1_co1_10), .S(
        early_found_msb_126_2_1_wmux_23_S), .Y(
        early_found_msb_126_2_1_y0_10), .FCO(
        early_found_msb_126_2_1_co0_11));
    CFG4 #( .INIT(16'h8CBF) )  \clkalign_curr_state_ns_5_0_.N_40_i  (
        .A(clkalign_curr_state_Z[3]), .B(clkalign_curr_state_Z[5]), .C(
        N_38), .D(N_25), .Y(N_40_i));
    SLE \early_late_end_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[1]));
    CFG3 #( .INIT(8'hD8) )  early_found_msb_127 (.A(emflag_cnt_Z[0]), 
        .B(N_2221), .C(N_2158), .Y(early_found_msb));
    SLE \tapcnt_final[5]  (.D(tapcnt_final_11[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_11_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(tapcnt_final_Z[5]));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_26 (.A(
        late_found_lsb_126_2_1_y0_11), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[51]), .D(late_flags_lsb_Z[115]), .FCI(
        late_found_lsb_126_2_1_co0_12), .S(
        late_found_lsb_126_2_1_wmux_26_S), .Y(
        late_found_lsb_126_2_1_y3_1), .FCO(
        late_found_lsb_126_2_1_co1_12));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_20 (.A(
        early_found_lsb_63_2_1_y0_9), .B(early_found_lsb_63_2_1_y3_0), 
        .C(early_found_lsb_63_2_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co0_9), .S(
        early_found_lsb_63_2_1_wmux_20_S), .Y(
        early_found_lsb_63_2_1_0_y21), .FCO(
        early_found_lsb_63_2_1_co1_9));
    CFG3 #( .INIT(8'h47) )  \clkalign_curr_state_ns_5_0_.m101  (.A(
        clkalign_curr_state_Z[0]), .B(clkalign_curr_state_Z[4]), .C(
        N_101), .Y(N_102));
    CFG4 #( .INIT(16'h7BDE) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state63_NE_2  (.A(
        tapcnt_final_Z[2]), .B(tapcnt_final_Z[1]), .C(tap_cnt_Z[2]), 
        .D(tap_cnt_Z[1]), .Y(clkalign_curr_state63_NE_2));
    SLE \late_flags_lsb[10]  (.D(late_flags_lsb_Z[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[10]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[4]), 
        .D(late_flags_lsb_Z[68]), .FCI(late_found_lsb_63_2_1_co1_4), 
        .S(late_found_lsb_63_2_1_wmux_11_S), .Y(
        late_found_lsb_63_2_1_y0_5), .FCO(late_found_lsb_63_2_1_co0_5));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNI5JTD3[3]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[3]), 
        .D(GND), .FCI(tapcnt_offset_cry[2]), .S(tapcnt_offset_s[3]), 
        .Y(tapcnt_offset_RNI5JTD3_Y[3]), .FCO(tapcnt_offset_cry[3]));
    SLE \late_flags_msb[125]  (.D(late_flags_msb_Z[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[125]));
    SLE \late_flags_msb[110]  (.D(late_flags_msb_Z[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[110]));
    SLE \late_flags_lsb[106]  (.D(late_flags_lsb_Z[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[106]));
    CFG4 #( .INIT(16'hFF40) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_6_0_0_933  
        (.A(rx_err_Z), .B(calc_done_Z), .C(clkalign_curr_state_Z[3]), 
        .D(un1_clkalign_curr_state_0_sqmuxa_6_0_0_933_1), .Y(N_2939));
    SLE \early_flags_lsb[26]  (.D(early_flags_lsb_Z[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[26]));
    CFG4 #( .INIT(16'h0F88) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state_1_sqmuxa_1_0_a3_RNIN2AC_0  
        (.A(N_643), .B(N_644), .C(tap_cnt_Z[7]), .D(
        clkalign_curr_state_1_sqmuxa_1), .Y(un1_early_flags_lsb14_1_i));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_24 (.A(
        late_found_lsb_126_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[35]), .D(late_flags_lsb_Z[99]), .FCI(
        late_found_lsb_126_2_1_co0_11), .S(
        late_found_lsb_126_2_1_wmux_24_S), .Y(
        late_found_lsb_126_2_1_y1_1), .FCO(
        late_found_lsb_126_2_1_co1_11));
    SLE \early_flags_lsb[104]  (.D(early_flags_lsb_Z[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[104]));
    SLE \late_flags_msb[56]  (.D(late_flags_msb_Z[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[56]));
    SLE \early_flags_lsb[68]  (.D(early_flags_lsb_Z[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[68]));
    CFG4 #( .INIT(16'hF1FF) )  
        \clkalign_curr_state_ns_5_0_.emflag_cnt10_i_0  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[4]), .C(
        clkalign_curr_state_Z[5]), .D(clkalign_curr_state_Z[0]), .Y(
        emflag_cnt10_i_0));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_41 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[30])
        , .D(late_flags_msb_Z[94]), .FCI(late_found_msb_63_2_1_co1_19), 
        .S(late_found_msb_63_2_1_wmux_41_S), .Y(
        late_found_msb_63_2_1_y0_18), .FCO(
        late_found_msb_63_2_1_co0_20));
    SLE \late_flags_msb[53]  (.D(late_flags_msb_Z[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[53]));
    CFG4 #( .INIT(16'hFFE0) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_0_sqmuxa_3_0  
        (.A(un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0), .B(
        un1_clkalign_curr_state_0_sqmuxa_3_0_a3_0_0), .C(N_125_mux), 
        .D(RX_RESET_LANE5), .Y(un1_clkalign_curr_state_0_sqmuxa_3_0));
    SLE late_not_found_lsb_d (.D(late_found_lsb_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(late_not_found_lsb_d_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_found_msb_63_2_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_msb_Z[8])
        , .D(early_flags_msb_Z[72]), .FCI(early_found_msb_63_2_1_co1_0)
        , .S(early_found_msb_63_2_1_wmux_3_S), .Y(
        early_found_msb_63_2_1_y0_1), .FCO(
        early_found_msb_63_2_1_co0_1));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNO[7]  (.A(VCC), .B(
        clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[7]), .D(
        GND), .FCI(tapcnt_offset_cry[6]), .S(tapcnt_offset_s[7]), .Y(
        tapcnt_offset_RNO_Y[7]), .FCO(tapcnt_offset_RNO_FCO[7]));
    SLE \early_flags_msb[9]  (.D(early_flags_msb_Z[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[9]));
    SLE \late_flags_lsb[91]  (.D(late_flags_lsb_Z[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[91]));
    CFG2 #( .INIT(4'h8) )  early_late_start_and_end_set5 (.A(
        early_late_end_set_Z), .B(early_late_start_set_Z), .Y(
        early_late_start_and_end_set5_Z));
    SLE \rst_cnt[5]  (.D(rst_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[5]));
    SLE \late_flags_msb[111]  (.D(late_flags_msb_Z[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[111]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_126_2_1_wmux_33 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        early_found_lsb_126_2_1_co1_15), .S(
        early_found_lsb_126_2_1_wmux_33_S), .Y(
        early_found_lsb_126_2_1_wmux_33_Y), .FCO(
        early_found_lsb_126_2_1_co0_16));
    SLE \tap_cnt[0]  (.D(tap_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tap_cnte), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tap_cnt_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_63_2_1_wmux_23 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[2]), 
        .D(late_flags_lsb_Z[66]), .FCI(late_found_lsb_63_2_1_co1_10), 
        .S(late_found_lsb_63_2_1_wmux_23_S), .Y(
        late_found_lsb_63_2_1_y0_10), .FCO(
        late_found_lsb_63_2_1_co0_11));
    SLE \early_flags_msb[65]  (.D(early_flags_msb_Z[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[65]));
    SLE \tapcnt_offset[5]  (.D(tapcnt_offset_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(tapcnt_offsete), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(tapcnt_offset_Z[5]));
    CFG4 #( .INIT(16'h0008) )  
        \clkalign_curr_state_ns_5_0_.early_late_start_set5_0_a3_1  (.A(
        clkalign_curr_state_Z[2]), .B(clkalign_curr_state_Z[0]), .C(
        N_533), .D(N_523), .Y(early_late_start_set5_0_a3_1));
    SLE \early_flags_msb[54]  (.D(early_flags_msb_Z[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[54]));
    SLE \early_late_end_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[0]));
    SLE \early_flags_lsb[28]  (.D(early_flags_lsb_Z[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[28]));
    SLE \early_flags_lsb[19]  (.D(early_flags_lsb_Z[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[19]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[7]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[7]), .D(early_late_init_val_Z[7]), .Y(
        tapcnt_final_11_iv_1[7]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_38 (.A(
        early_found_msb_126_2_1_y0_16), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[55]), .D(early_flags_msb_Z[119]), .FCI(
        early_found_msb_126_2_1_co0_18), .S(
        early_found_msb_126_2_1_wmux_38_S), .Y(
        early_found_msb_126_2_1_y3_2), .FCO(
        early_found_msb_126_2_1_co1_18));
    CFG4 #( .INIT(16'h2075) )  \clkalign_curr_state_ns_5_0_.m76  (.A(
        clkalign_curr_state_Z[5]), .B(clkalign_curr_state_Z[3]), .C(
        N_75), .D(N_71), .Y(clkalign_curr_state_ns[1]));
    SLE \sig_tapcnt_final_2[7]  (.D(un2_sig_tapcnt_final_2_cry_7_Z), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[7]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_126_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[21])
        , .D(late_flags_msb_Z[85]), .FCI(late_found_msb_126_2_1_co1_5), 
        .S(late_found_msb_126_2_1_wmux_13_S), .Y(
        late_found_msb_126_2_1_y0_6), .FCO(
        late_found_msb_126_2_1_co0_6));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_0 (.A(
        early_found_msb_126_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[33]), .D(early_flags_msb_Z[97]), .FCI(
        early_found_msb_126_2_1_0_co0), .S(
        early_found_msb_126_2_1_wmux_0_S), .Y(
        early_found_msb_126_2_1_0_y1), .FCO(
        early_found_msb_126_2_1_0_co1));
    SLE \late_flags_lsb[95]  (.D(late_flags_lsb_Z[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[95]));
    ARI1 #( .INIT(20'h0CEC2) )  early_found_lsb_63_2_1_wmux_10 (.A(
        early_found_lsb_63_2_1_0_y21), .B(early_found_lsb_63_2_1_0_y9), 
        .C(emflag_cnt_Z[2]), .D(emflag_cnt_Z[1]), .FCI(
        early_found_lsb_63_2_1_co0_4), .S(
        early_found_lsb_63_2_1_wmux_10_S), .Y(
        early_found_lsb_63_2_1_y0_4), .FCO(
        early_found_lsb_63_2_1_co1_4));
    SLE \late_flags_lsb[57]  (.D(late_flags_lsb_Z[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[57]));
    ARI1 #( .INIT(20'h48800) )  \tapcnt_offset_RNIADF02[1]  (.A(VCC), 
        .B(clkalign_curr_state_RNIJB1J_Y[0]), .C(tapcnt_offset_Z[1]), 
        .D(GND), .FCI(tapcnt_offset_cry[0]), .S(tapcnt_offset_s[1]), 
        .Y(tapcnt_offset_RNIADF02_Y[1]), .FCO(tapcnt_offset_cry[1]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_126_2_1_wmux_19 (.A(
        late_found_msb_126_2_1_y7_0), .B(late_found_msb_126_2_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co1_8), .S(
        late_found_msb_126_2_1_wmux_19_S), .Y(
        late_found_msb_126_2_1_y0_9), .FCO(
        late_found_msb_126_2_1_co0_9));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_1 (.A(
        early_late_init_val_Z[1]), .B(early_late_nxt_val_Z[1]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_0_Z), .S(
        un2_sig_tapcnt_final_2_cry_1_S), .Y(
        un2_sig_tapcnt_final_2_cry_1_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_1_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_126_2_1_wmux_31 (.A(
        early_found_lsb_126_2_1_y7_1), .B(early_found_lsb_126_2_1_y5_1)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_126_2_1_co1_14), .S(
        early_found_lsb_126_2_1_wmux_31_S), .Y(
        early_found_lsb_126_2_1_y0_14), .FCO(
        early_found_lsb_126_2_1_co0_15));
    CFG4 #( .INIT(16'h193B) )  \clkalign_curr_state_ns_5_0_.m37_2_1_1  
        (.A(clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), 
        .C(N_134_mux), .D(N_30), .Y(m37_2_1_1));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_6 (.A(
        early_late_init_val_Z[6]), .B(early_late_nxt_val_Z[6]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_5_Z), .S(
        un2_sig_tapcnt_final_2_cry_6_S), .Y(
        un2_sig_tapcnt_final_2_cry_6_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_6_Z));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_2 
        (.A(early_late_nxt_val_Z[2]), .B(early_late_init_val_Z[2]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_1_Z), 
        .S(early_late_init_nxt_val_status5_cry_2_S), .Y(
        early_late_init_nxt_val_status5_cry_2_Y), .FCO(
        early_late_init_nxt_val_status5_cry_2_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_126_2_1_wmux_35 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_lsb_Z[7])
        , .D(early_flags_lsb_Z[71]), .FCI(
        early_found_lsb_126_2_1_co1_16), .S(
        early_found_lsb_126_2_1_wmux_35_S), .Y(
        early_found_lsb_126_2_1_y0_15), .FCO(
        early_found_lsb_126_2_1_co0_17));
    SLE \sig_tapcnt_final_2[1]  (.D(sig_tapcnt_final_2_3_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[1]));
    SLE \late_flags_msb[12]  (.D(late_flags_msb_Z[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[12]));
    SLE start_trng_fg (.D(start_trng_fg6), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(start_trng_fg_Z));
    SLE \early_flags_msb[51]  (.D(early_flags_msb_Z[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[51]));
    SLE \early_flags_lsb[59]  (.D(early_flags_lsb_Z[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[59]));
    ARI1 #( .INIT(20'h555AA) )  un2_sig_tapcnt_final_2_cry_3 (.A(
        early_late_init_val_Z[3]), .B(early_late_nxt_val_Z[3]), .C(GND)
        , .D(GND), .FCI(un2_sig_tapcnt_final_2_cry_2_Z), .S(
        un2_sig_tapcnt_final_2_cry_3_S), .Y(
        un2_sig_tapcnt_final_2_cry_3_Y), .FCO(
        un2_sig_tapcnt_final_2_cry_3_Z));
    SLE \early_late_start_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[6]));
    SLE \early_flags_lsb[80]  (.D(early_flags_lsb_Z[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[80]));
    CFG4 #( .INIT(16'h0001) )  
        \clkalign_curr_state_ns_5_0_.un1_early_late_end_set12_3_i_0_RNI81D21  
        (.A(clkalign_curr_state_Z[5]), .B(
        un1_early_late_end_set12_3_i_0), .C(N_525), .D(N_619), .Y(
        N_515_i));
    SLE early_found_lsb_d (.D(early_found_lsb), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(early_found_lsb_d_Z));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_msb_126_2_1_wmux_44 (.A(
        early_found_msb_126_2_1_y0_19), .B(
        early_found_msb_126_2_1_y3_2), .C(early_found_msb_126_2_1_y1_2)
        , .D(emflag_cnt_Z[3]), .FCI(early_found_msb_126_2_1_co0_21), 
        .S(early_found_msb_126_2_1_wmux_44_S), .Y(
        early_found_msb_126_2_1_0_y45), .FCO(
        early_found_msb_126_2_1_co1_21));
    SLE \early_flags_lsb[73]  (.D(early_flags_lsb_Z[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[73]));
    ARI1 #( .INIT(20'h48800) )  \tap_cnt_cry[2]  (.A(VCC), .B(
        tap_cnt_cry_cy_Y[0]), .C(tap_cnt_Z[2]), .D(GND), .FCI(
        tap_cnt_cry_Z[1]), .S(tap_cnt_s[2]), .Y(tap_cnt_cry_Y[2]), 
        .FCO(tap_cnt_cry_Z[2]));
    SLE \early_flags_msb[56]  (.D(early_flags_msb_Z[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[56]));
    SLE \late_flags_msb[115]  (.D(late_flags_msb_Z[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[115]));
    CFG2 #( .INIT(4'h6) )  \clkalign_curr_state_ns_5_0_.SUM_0_0_x2[1]  
        (.A(CO0_0), .B(cnt_Z[1]), .Y(N_554_i));
    SLE \early_late_end_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_late_end_set12_1_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_end_val_Z[6]));
    CFG2 #( .INIT(4'h4) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_0_sqmuxa_1  (.A(
        N_538_i), .B(clkalign_curr_state_d[27]), .Y(
        tapcnt_final_0_sqmuxa_1));
    ARI1 #( .INIT(20'h0FA44) )  early_found_lsb_63_2_1_wmux_29 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[26]), .D(early_flags_lsb_Z[90]), .FCI(
        early_found_lsb_63_2_1_co1_13), .S(
        early_found_lsb_63_2_1_wmux_29_S), .Y(
        early_found_lsb_63_2_1_y0_13), .FCO(
        early_found_lsb_63_2_1_co0_14));
    SLE \sig_tapcnt_final_2[3]  (.D(sig_tapcnt_final_2_3_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(sig_tapcnt_final_2_Z[3]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_30 (.A(
        early_found_msb_126_2_1_y0_13), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[59]), .D(early_flags_msb_Z[123]), .FCI(
        early_found_msb_126_2_1_co0_14), .S(
        early_found_msb_126_2_1_wmux_30_S), .Y(
        early_found_msb_126_2_1_y7_1), .FCO(
        early_found_msb_126_2_1_co1_14));
    SLE \clkalign_curr_state[3]  (.D(clkalign_curr_state_ns[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(clkalign_curr_state_Z[3]));
    SLE \late_flags_lsb[102]  (.D(late_flags_lsb_Z[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[102]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_msb_126_2_1_wmux_8 (.A(
        late_found_msb_126_2_1_y0_3), .B(late_found_msb_126_2_1_0_y3), 
        .C(late_found_msb_126_2_1_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co0_3), .S(
        late_found_msb_126_2_1_wmux_8_S), .Y(
        late_found_msb_126_2_1_0_y9), .FCO(
        late_found_msb_126_2_1_co1_3));
    SLE \late_flags_lsb[54]  (.D(late_flags_lsb_Z[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[54]));
    SLE \early_late_init_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[1]));
    SLE \late_flags_lsb[68]  (.D(late_flags_lsb_Z[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[68]));
    SLE \early_flags_lsb[117]  (.D(early_flags_lsb_Z[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[117]));
    CFG4 #( .INIT(16'h5111) )  \clkalign_curr_state_ns_5_0_.m65  (.A(
        clkalign_curr_state_Z[1]), .B(N_19_i), .C(rx_err_Z), .D(
        calc_done_Z), .Y(i22_mux));
    SLE \early_flags_msb[117]  (.D(early_flags_msb_Z[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[117]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_s[7]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y[0]), .C(emflag_cnt_Z[7]), .D(GND), .FCI(
        emflag_cnt_cry_Z[6]), .S(emflag_cnt_s_Z[7]), .Y(
        emflag_cnt_s_Y[7]), .FCO(emflag_cnt_s_FCO[7]));
    CFG2 #( .INIT(4'h1) )  sig_tapcnt_final_111_3 (.A(
        early_late_end_val_Z[0]), .B(early_late_end_val_Z[3]), .Y(
        sig_tapcnt_final_111_3_Z));
    SLE \late_flags_msb[124]  (.D(late_flags_msb_Z[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[124]));
    CFG4 #( .INIT(16'hC480) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv_1[5]  (.A(
        early_late_init_nxt_val_status_Z), .B(tapcnt_final_2_sqmuxa_1), 
        .C(sig_tapcnt_final_2_Z[5]), .D(early_late_init_val_Z[5]), .Y(
        tapcnt_final_11_iv_1[5]));
    SLE \late_flags_lsb[40]  (.D(late_flags_lsb_Z[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[40]));
    SLE \early_flags_msb[58]  (.D(early_flags_msb_Z[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[58]));
    CFG4 #( .INIT(16'h0010) )  
        \clkalign_curr_state_ns_5_0_.un1_clkalign_curr_state_1_0_a3_0  
        (.A(clkalign_curr_state_Z[0]), .B(clkalign_curr_state_Z[2]), 
        .C(clkalign_curr_state_Z[4]), .D(clkalign_curr_state_Z[1]), .Y(
        un1_clkalign_curr_state_1_0_a3_0));
    CFG3 #( .INIT(8'hD8) )  late_found_msb_127 (.A(emflag_cnt_Z[0]), 
        .B(N_2348), .C(N_2285), .Y(late_found_msb));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_16 (.A(
        late_found_lsb_126_2_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[45]), .D(late_flags_lsb_Z[109]), .FCI(
        late_found_lsb_126_2_1_co0_7), .S(
        late_found_lsb_126_2_1_wmux_16_S), .Y(
        late_found_lsb_126_2_1_y5_0), .FCO(
        late_found_lsb_126_2_1_co1_7));
    SLE \late_flags_msb[48]  (.D(late_flags_msb_Z[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[48]));
    SLE \late_flags_lsb[26]  (.D(late_flags_lsb_Z[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[26]));
    SLE \early_flags_lsb[5]  (.D(early_flags_lsb_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[5]));
    SLE \late_flags_lsb[23]  (.D(late_flags_lsb_Z[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[23]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_0 
        (.A(early_late_nxt_val_Z[0]), .B(early_late_init_val_Z[0]), .C(
        GND), .D(GND), .FCI(GND), .S(
        early_late_init_nxt_val_status5_cry_0_S), .Y(
        early_late_init_nxt_val_status5_cry_0_Y), .FCO(
        early_late_init_nxt_val_status5_cry_0_Z));
    SLE late_not_found_msb_d (.D(late_found_msb_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(late_not_found_msb_d_Z));
    SLE \early_flags_msb[124]  (.D(early_flags_msb_Z[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[124]));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_63_2_1_wmux_36 (.A(
        late_found_msb_63_2_1_y0_15), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[38]), .D(late_flags_msb_Z[102]), .FCI(
        late_found_msb_63_2_1_co0_17), .S(
        late_found_msb_63_2_1_wmux_36_S), .Y(
        late_found_msb_63_2_1_y1_2), .FCO(late_found_msb_63_2_1_co1_17)
        );
    CFG4 #( .INIT(16'h8B03) )  
        \clkalign_curr_state_ns_5_0_.clkalign_curr_state63_NE_i_RNIJNDO2  
        (.A(clkalign_curr_state63), .B(clkalign_curr_state_Z[1]), .C(
        N_128_mux), .D(m44_0), .Y(N_46));
    CFG4 #( .INIT(16'h269D) )  \clkalign_curr_state_ns_5_0_.m23  (.A(
        clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[2]), .C(
        N_139_mux), .D(clkalign_curr_state_Z[4]), .Y(N_3109_mux));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_14 (.A(
        late_found_lsb_126_2_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[53]), .D(late_flags_lsb_Z[117]), .FCI(
        late_found_lsb_126_2_1_co0_6), .S(
        late_found_lsb_126_2_1_wmux_14_S), .Y(
        late_found_lsb_126_2_1_y3_0), .FCO(
        late_found_lsb_126_2_1_co1_6));
    SLE \early_late_init_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_14_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_init_val_Z[0]));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_lsb_63_2_1_wmux_19 (.A(
        early_found_lsb_63_2_1_y7_0), .B(early_found_lsb_63_2_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co1_8), .S(
        early_found_lsb_63_2_1_wmux_19_S), .Y(
        early_found_lsb_63_2_1_y0_9), .FCO(
        early_found_lsb_63_2_1_co0_9));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[3]  (.A(VCC), .B(
        rst_cnt_Z[3]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[2]), .S(
        rst_cnt_s[3]), .Y(rst_cnt_cry_Y[3]), .FCO(rst_cnt_cry_Z[3]));
    SLE \early_flags_msb[1]  (.D(early_flags_msb_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[1]));
    SLE \late_flags_lsb[86]  (.D(late_flags_lsb_Z[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[86]));
    ARI1 #( .INIT(20'h0FA0C) )  early_found_lsb_63_2_1_wmux_32 (.A(
        early_found_lsb_63_2_1_y0_14), .B(early_found_lsb_63_2_1_y3_1), 
        .C(early_found_lsb_63_2_1_y1_1), .D(emflag_cnt_Z[3]), .FCI(
        early_found_lsb_63_2_1_co0_15), .S(
        early_found_lsb_63_2_1_wmux_32_S), .Y(
        early_found_lsb_63_2_1_0_y33), .FCO(
        early_found_lsb_63_2_1_co1_15));
    SLE \late_flags_lsb[83]  (.D(late_flags_lsb_Z[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[83]));
    SLE \late_flags_msb[38]  (.D(late_flags_msb_Z[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[38]));
    SLE \clkalign_curr_state[4]  (.D(clkalign_curr_state_ns[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(clkalign_curr_state_Z[4]));
    SLE \rst_cnt[9]  (.D(rst_cnt_s_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        current_state_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(rst_cnt_Z[9]));
    CFG4 #( .INIT(16'h0001) )  clkalign_curr_state81_NE_i (.A(
        tapcnt_offset_Z[2]), .B(tapcnt_offset_Z[5]), .C(
        clkalign_curr_state81_NE_4_Z), .D(clkalign_curr_state81_NE_3_Z)
        , .Y(clkalign_curr_state81));
    ARI1 #( .INIT(20'h0F588) )  late_found_lsb_126_2_1_wmux_42 (.A(
        late_found_lsb_126_2_1_y0_18), .B(emflag_cnt_Z[5]), .C(
        late_flags_lsb_Z[63]), .D(late_flags_lsb_Z[127]), .FCI(
        late_found_lsb_126_2_1_co0_20), .S(
        late_found_lsb_126_2_1_wmux_42_S), .Y(
        late_found_lsb_126_2_1_y7_2), .FCO(
        late_found_lsb_126_2_1_co1_20));
    SLE \late_flags_lsb[30]  (.D(late_flags_lsb_Z[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[30]));
    SLE \early_flags_lsb[93]  (.D(early_flags_lsb_Z[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[93]));
    CFG4 #( .INIT(16'hDC76) )  \clkalign_curr_state_ns_5_0_.m16_2_0  (
        .A(clkalign_curr_state_Z[1]), .B(clkalign_curr_state_Z[4]), .C(
        N_12), .D(m16_2_0_1_0), .Y(m16_2_0));
    ARI1 #( .INIT(20'h4AA00) )  rst_cnt_s_1133 (.A(VCC), .B(
        rst_cnt_Z[0]), .C(GND), .D(GND), .FCI(VCC), .S(
        rst_cnt_s_1133_S), .Y(rst_cnt_s_1133_Y), .FCO(
        rst_cnt_s_1133_FCO));
    SLE \early_late_start_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[2]));
    SLE \early_flags_msb[104]  (.D(early_flags_msb_Z[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[104]));
    ARI1 #( .INIT(20'h0F588) )  early_found_msb_126_2_1_wmux_24 (.A(
        early_found_msb_126_2_1_y0_10), .B(emflag_cnt_Z[5]), .C(
        early_flags_msb_Z[35]), .D(early_flags_msb_Z[99]), .FCI(
        early_found_msb_126_2_1_co0_11), .S(
        early_found_msb_126_2_1_wmux_24_S), .Y(
        early_found_msb_126_2_1_y1_1), .FCO(
        early_found_msb_126_2_1_co1_11));
    SLE \late_flags_msb[88]  (.D(late_flags_msb_Z[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[88]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_init_nxt_val_status5_cry_7 
        (.A(early_late_nxt_val_Z[7]), .B(early_late_init_val_Z[7]), .C(
        GND), .D(GND), .FCI(early_late_init_nxt_val_status5_cry_6_Z), 
        .S(early_late_init_nxt_val_status5_cry_7_S), .Y(
        early_late_init_nxt_val_status5_cry_7_Y), .FCO(
        early_late_init_nxt_val_status5));
    ARI1 #( .INIT(20'h0F588) )  late_found_msb_126_2_1_wmux_0 (.A(
        late_found_msb_126_2_1_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_msb_Z[33]), .D(late_flags_msb_Z[97]), .FCI(
        late_found_msb_126_2_1_0_co0), .S(
        late_found_msb_126_2_1_wmux_0_S), .Y(
        late_found_msb_126_2_1_0_y1), .FCO(
        late_found_msb_126_2_1_0_co1));
    ARI1 #( .INIT(20'h0F588) )  early_found_lsb_126_2_1_wmux_40 (.A(
        early_found_lsb_126_2_1_y0_17), .B(emflag_cnt_Z[5]), .C(
        early_flags_lsb_Z[47]), .D(early_flags_lsb_Z[111]), .FCI(
        early_found_lsb_126_2_1_co0_19), .S(
        early_found_lsb_126_2_1_wmux_40_S), .Y(
        early_found_lsb_126_2_1_y5_2), .FCO(
        early_found_lsb_126_2_1_co1_19));
    ARI1 #( .INIT(20'h42200) )  \clkalign_curr_state_RNIJB1J[0]  (.A(
        VCC), .B(clkalign_curr_state_Z[0]), .C(
        clkalign_curr_state_Z[3]), .D(GND), .FCI(VCC), .S(
        clkalign_curr_state_RNIJB1J_S[0]), .Y(
        clkalign_curr_state_RNIJB1J_Y[0]), .FCO(tapcnt_offset_cry_cy));
    SLE \late_flags_msb[66]  (.D(late_flags_msb_Z[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[66]));
    CFG2 #( .INIT(4'hE) )  
        \clkalign_curr_state_ns_5_0_.tapcnt_final_11_iv[7]  (.A(
        tapcnt_final_11_iv_1[7]), .B(tapcnt_final_11_iv_0[7]), .Y(
        tapcnt_final_11[7]));
    SLE \early_flags_msb[47]  (.D(early_flags_msb_Z[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[47]));
    SLE \late_flags_msb[63]  (.D(late_flags_msb_Z[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[63]));
    SLE \early_flags_msb[83]  (.D(early_flags_msb_Z[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[83]));
    SLE \early_flags_lsb[62]  (.D(early_flags_lsb_Z[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[62]));
    ARI1 #( .INIT(20'h0FA44) )  late_found_lsb_126_2_1_wmux_27 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_lsb_Z[11])
        , .D(late_flags_lsb_Z[75]), .FCI(late_found_lsb_126_2_1_co1_12)
        , .S(late_found_lsb_126_2_1_wmux_27_S), .Y(
        late_found_lsb_126_2_1_y0_12), .FCO(
        late_found_lsb_126_2_1_co0_13));
    SLE \late_flags_msb[114]  (.D(late_flags_msb_Z[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[114]));
    SLE \early_late_start_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_clkalign_curr_state_15_0), .ALn(current_state_0), .ADn(VCC)
        , .SLn(N_677_i), .SD(GND), .LAT(GND), .Q(
        early_late_start_val_Z[0]));
    SLE \early_flags_lsb[33]  (.D(early_flags_lsb_Z[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[33]));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_63_2_1_wmux_21 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_63_2_1_co1_9), .S(
        late_found_lsb_63_2_1_wmux_21_S), .Y(
        late_found_lsb_63_2_1_wmux_21_Y), .FCO(
        late_found_lsb_63_2_1_co0_10));
    ARI1 #( .INIT(20'h0FA0C) )  late_found_lsb_126_2_1_wmux_22 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[4]), .D(VCC), .FCI(
        late_found_lsb_126_2_1_co0_10), .S(
        late_found_lsb_126_2_1_wmux_22_S), .Y(
        late_found_lsb_126_2_1_wmux_22_Y), .FCO(
        late_found_lsb_126_2_1_co1_10));
    SLE \late_flags_msb[17]  (.D(late_flags_msb_Z[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[17]));
    SLE \early_flags_msb[3]  (.D(early_flags_msb_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[3]));
    SLE \early_flags_msb[23]  (.D(early_flags_msb_Z[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[23]));
    SLE \late_flags_msb[72]  (.D(late_flags_msb_Z[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[72]));
    SLE \early_flags_msb[19]  (.D(early_flags_msb_Z[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[19]));
    ARI1 #( .INIT(20'h5AA55) )  early_late_start_end_val_status5_cry_1 
        (.A(early_late_end_val_Z[1]), .B(early_late_start_val_Z[1]), 
        .C(GND), .D(GND), .FCI(
        early_late_start_end_val_status5_cry_0_Z), .S(
        early_late_start_end_val_status5_cry_1_S), .Y(
        early_late_start_end_val_status5_cry_1_Y), .FCO(
        early_late_start_end_val_status5_cry_1_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_found_msb_126_2_1_wmux_19 (.A(
        early_found_msb_126_2_1_y7_0), .B(early_found_msb_126_2_1_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_found_msb_126_2_1_co1_8), .S(
        early_found_msb_126_2_1_wmux_19_S), .Y(
        early_found_msb_126_2_1_y0_9), .FCO(
        early_found_msb_126_2_1_co0_9));
    SLE \late_flags_lsb[69]  (.D(late_flags_lsb_Z[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(late_flags_lsb_Z[69]));
    SLE \early_flags_msb[123]  (.D(early_flags_msb_Z[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(early_flags_msb_Z[123]));
    SLE \early_flags_lsb[4]  (.D(early_flags_lsb_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[4]));
    SLE \early_flags_lsb[22]  (.D(early_flags_lsb_Z[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        un1_early_flags_lsb14_1_i), .ALn(current_state_0), .ADn(VCC), 
        .SLn(N_673_i), .SD(GND), .LAT(GND), .Q(early_flags_lsb_Z[22]));
    ARI1 #( .INIT(20'h0EC2C) )  late_found_msb_126_2_1_wmux_31 (.A(
        late_found_msb_126_2_1_y7_1), .B(late_found_msb_126_2_1_y5_1), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_found_msb_126_2_1_co1_14), .S(
        late_found_msb_126_2_1_wmux_31_S), .Y(
        late_found_msb_126_2_1_y0_14), .FCO(
        late_found_msb_126_2_1_co0_15));
    ARI1 #( .INIT(20'h0FA44) )  late_found_msb_63_2_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_msb_Z[20])
        , .D(late_flags_msb_Z[84]), .FCI(late_found_msb_63_2_1_co1_5), 
        .S(late_found_msb_63_2_1_wmux_13_S), .Y(
        late_found_msb_63_2_1_y0_6), .FCO(late_found_msb_63_2_1_co0_6));
    SLE \late_flags_msb[49]  (.D(late_flags_msb_Z[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_early_flags_lsb14_i), 
        .ALn(current_state_0), .ADn(VCC), .SLn(N_673_i), .SD(GND), 
        .LAT(GND), .Q(late_flags_msb_Z[49]));
    CFG3 #( .INIT(8'h47) )  \clkalign_curr_state_ns_5_0_.m16_2_0_1_0  
        (.A(clkalign_curr_state_Z[0]), .B(clkalign_curr_state_Z[4]), 
        .C(N_5), .Y(m16_2_0_1_0));
    
endmodule


module 
        PF_IOD_GENERIC_RX_C1_TR_PF_IOD_GENERIC_RX_C1_TR_0_COREBCLKSCLKALIGN_Z2(
        
       current_state_0,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV,
       COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE,
       CLK_TRAIN_ERROR_c,
       PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE,
       PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE
    );
input  current_state_0;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
output RX_CLK_ALIGN_DONE_arst;
input  PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0;
input  PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV;
output COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE;
output CLK_TRAIN_ERROR_c;
output PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE;
input  PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE;

    wire GND, VCC;
    
    ICB_BCLKSCLKALIGN_Z3 \genblk1.U_ICB_BCLKSCLKALIGN  (
        .current_state_0(current_state_0), 
        .PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), 
        .PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE(
        PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE), .CLK_TRAIN_ERROR_c(
        CLK_TRAIN_ERROR_c), .COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE(
        COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), 
        .RX_CLK_ALIGN_DONE_arst(RX_CLK_ALIGN_DONE_arst), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1_TR(
       current_state_0,
       PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE,
       PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE,
       CLK_TRAIN_ERROR_c,
       COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD,
       COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0,
       PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0,
       RX_CLK_ALIGN_DONE_arst,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G
    );
input  current_state_0;
input  PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE;
output PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE;
output CLK_TRAIN_ERROR_c;
output COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD;
output COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS;
input  PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0;
input  PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0;
output RX_CLK_ALIGN_DONE_arst;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;

    wire GND, VCC;
    
    
        PF_IOD_GENERIC_RX_C1_TR_PF_IOD_GENERIC_RX_C1_TR_0_COREBCLKSCLKALIGN_Z2 
        PF_IOD_GENERIC_RX_C1_TR_0 (.current_state_0(current_state_0), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV), 
        .COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE(
        COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE), .CLK_TRAIN_ERROR_c(
        CLK_TRAIN_ERROR_c), .PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE(
        PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE), 
        .PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_RX_C1(
       BIT_ALGN_EYE_IN_c,
       RXD_N,
       RXD,
       rev_bits_0_out_data_4,
       EYE_MONITOR_EARLY_net_0,
       EYE_MONITOR_LATE_net_0,
       ACT_UNIQUE_rev_bits_0_out_data,
       current_state_0,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD,
       BIT_ALGN_OOR_0_c,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD,
       BIT_ALGN_OOR_c,
       RX_CLK_ALIGN_DONE_arst,
       CLK_TRAIN_ERROR_c,
       RX_CLK_P,
       RX_CLK_N,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G
    );
input  [2:0] BIT_ALGN_EYE_IN_c;
input  [1:0] RXD_N;
input  [1:0] RXD;
output [7:0] rev_bits_0_out_data_4;
output [1:0] EYE_MONITOR_EARLY_net_0;
output [1:0] EYE_MONITOR_LATE_net_0;
output [7:0] ACT_UNIQUE_rev_bits_0_out_data;
input  current_state_0;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR;
input  CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD;
output BIT_ALGN_OOR_0_c;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR;
input  CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD;
output BIT_ALGN_OOR_c;
output RX_CLK_ALIGN_DONE_arst;
output CLK_TRAIN_ERROR_c;
input  RX_CLK_P;
input  RX_CLK_N;
output PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;

    wire [2:0] PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT;
    wire [2:0] PF_LANECTRL_0_FIFO_RD_PTR;
    wire [2:0] PF_LANECTRL_0_FIFO_WR_PTR;
    wire [0:0] PF_LANECTRL_0_RX_DQS_90;
    wire HS_IO_CLK_CASCADED_Y, Y_0, HS_IO_CLK_FIFO_Y, Y_1, 
        PF_CLK_DIV_FIFO_CLK_DIV_OUT, CLK_0_Y, PAUSE_MX_0_Y, 
        COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE, GND, 
        PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE, 
        PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK, HS_IO_CLK_RX_Y, 
        PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK, 
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE, 
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV, 
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD, 
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS, 
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0, 
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0, 
        PF_LANECTRL_0_TX_SYNC_RST, PF_LANECTRL_0_RX_SYNC_RST, 
        PF_LANECTRL_0_ARST_N, VCC;
    
    PF_IOD_GENERIC_RX_C1_PF_CLK_DIV_RXCLK_PF_CLK_DIV_DELAY 
        PF_CLK_DIV_RXCLK (.PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK(
        PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK), .HS_IO_CLK_CASCADED_Y(
        HS_IO_CLK_CASCADED_Y));
    CLKINT CLKINT_0 (.A(PF_CLK_DIV_FIFO_CLK_DIV_OUT), .Y(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G));
    CLKINT HS_IO_CLK_CASCADED_RNIIIH5 (.A(Y_0), .Y(
        HS_IO_CLK_CASCADED_Y));
    INBUF_DIFF CLK_0 (.PADP(RX_CLK_P), .PADN(RX_CLK_N), .Y(CLK_0_Y));
    PF_IOD_GENERIC_RX_C1_PF_CLK_DIV_FIFO_PF_CLK_DIV_DELAY 
        PF_CLK_DIV_FIFO (.PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK(
        PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK), 
        .PF_CLK_DIV_FIFO_CLK_DIV_OUT(PF_CLK_DIV_FIFO_CLK_DIV_OUT), 
        .HS_IO_CLK_CASCADED_Y(HS_IO_CLK_CASCADED_Y), 
        .PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV));
    HS_IO_CLK HS_IO_CLK_RX (.A(PF_CLK_DIV_RXCLK_CLK_OUT_HS_IO_CLK), .Y(
        HS_IO_CLK_RX_Y));
    HS_IO_CLK HS_IO_CLK_FIFO (.A(PF_CLK_DIV_FIFO_CLK_OUT_HS_IO_CLK), 
        .Y(Y_1));
    GND GND_Z (.Y(GND));
    PF_IOD_GENERIC_RX_C1_PF_IOD_CLK_TRAINING_PF_IOD 
        PF_IOD_CLK_TRAINING (.PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), .HS_IO_CLK_FIFO_Y(
        HS_IO_CLK_FIFO_Y), .PF_LANECTRL_0_TX_SYNC_RST(
        PF_LANECTRL_0_TX_SYNC_RST), .PF_LANECTRL_0_RX_SYNC_RST(
        PF_LANECTRL_0_RX_SYNC_RST), .PF_LANECTRL_0_ARST_N(
        PF_LANECTRL_0_ARST_N), .PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS));
    CLKINT HS_IO_CLK_FIFO_RNIEMED (.A(Y_1), .Y(HS_IO_CLK_FIFO_Y));
    HS_IO_CLK HS_IO_CLK_CASCADED (.A(CLK_0_Y), .Y(Y_0));
    PF_IOD_GENERIC_RX_C1_PF_LANECTRL_0_PF_LANECTRL PF_LANECTRL_0 (
        .PF_LANECTRL_0_FIFO_RD_PTR({PF_LANECTRL_0_FIFO_RD_PTR[2], 
        PF_LANECTRL_0_FIFO_RD_PTR[1], PF_LANECTRL_0_FIFO_RD_PTR[0]}), 
        .PF_LANECTRL_0_FIFO_WR_PTR({PF_LANECTRL_0_FIFO_WR_PTR[2], 
        PF_LANECTRL_0_FIFO_WR_PTR[1], PF_LANECTRL_0_FIFO_WR_PTR[0]}), 
        .PF_LANECTRL_0_RX_DQS_90_0(PF_LANECTRL_0_RX_DQS_90[0]), 
        .PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), .BIT_ALGN_EYE_IN_c({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .current_state_0(current_state_0), 
        .PAUSE_MX_0_Y(PAUSE_MX_0_Y), .PF_LANECTRL_0_TX_SYNC_RST(
        PF_LANECTRL_0_TX_SYNC_RST), .PF_LANECTRL_0_RX_SYNC_RST(
        PF_LANECTRL_0_RX_SYNC_RST), .PF_LANECTRL_0_ARST_N(
        PF_LANECTRL_0_ARST_N), .HS_IO_CLK_RX_Y(HS_IO_CLK_RX_Y), 
        .HS_IO_CLK_FIFO_Y(HS_IO_CLK_FIFO_Y), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G));
    PF_IOD_GENERIC_RX_C1_PF_IOD_RX_PF_IOD PF_IOD_RX (
        .ACT_UNIQUE_rev_bits_0_out_data({
        ACT_UNIQUE_rev_bits_0_out_data[7], 
        ACT_UNIQUE_rev_bits_0_out_data[6], 
        ACT_UNIQUE_rev_bits_0_out_data[5], 
        ACT_UNIQUE_rev_bits_0_out_data[4], 
        ACT_UNIQUE_rev_bits_0_out_data[3], 
        ACT_UNIQUE_rev_bits_0_out_data[2], 
        ACT_UNIQUE_rev_bits_0_out_data[1], 
        ACT_UNIQUE_rev_bits_0_out_data[0]}), .EYE_MONITOR_LATE_net_0({
        EYE_MONITOR_LATE_net_0[1], EYE_MONITOR_LATE_net_0[0]}), 
        .EYE_MONITOR_EARLY_net_0({EYE_MONITOR_EARLY_net_0[1], 
        EYE_MONITOR_EARLY_net_0[0]}), 
        .PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT({
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[2], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[1], 
        PF_LANECTRL_0_EYE_MONITOR_WIDTH_OUT[0]}), 
        .PF_LANECTRL_0_FIFO_RD_PTR({PF_LANECTRL_0_FIFO_RD_PTR[2], 
        PF_LANECTRL_0_FIFO_RD_PTR[1], PF_LANECTRL_0_FIFO_RD_PTR[0]}), 
        .PF_LANECTRL_0_FIFO_WR_PTR({PF_LANECTRL_0_FIFO_WR_PTR[2], 
        PF_LANECTRL_0_FIFO_WR_PTR[1], PF_LANECTRL_0_FIFO_WR_PTR[0]}), 
        .PF_LANECTRL_0_RX_DQS_90_0(PF_LANECTRL_0_RX_DQS_90[0]), 
        .rev_bits_0_out_data_4({rev_bits_0_out_data_4[7], 
        rev_bits_0_out_data_4[6], rev_bits_0_out_data_4[5], 
        rev_bits_0_out_data_4[4], rev_bits_0_out_data_4[3], 
        rev_bits_0_out_data_4[2], rev_bits_0_out_data_4[1], 
        rev_bits_0_out_data_4[0]}), .RXD({RXD[1], RXD[0]}), .RXD_N({
        RXD_N[1], RXD_N[0]}), .BIT_ALGN_OOR_c(BIT_ALGN_OOR_c), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS), .HS_IO_CLK_FIFO_Y(
        HS_IO_CLK_FIFO_Y), .PF_LANECTRL_0_TX_SYNC_RST(
        PF_LANECTRL_0_TX_SYNC_RST), .PF_LANECTRL_0_RX_SYNC_RST(
        PF_LANECTRL_0_RX_SYNC_RST), .PF_LANECTRL_0_ARST_N(
        PF_LANECTRL_0_ARST_N), .BIT_ALGN_OOR_0_c(BIT_ALGN_OOR_0_c), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS));
    VCC VCC_Z (.Y(VCC));
    MX2 PAUSE_MX_0 (.A(COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE), .B(
        GND), .S(PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE), .Y(
        PAUSE_MX_0_Y));
    PF_IOD_GENERIC_RX_C1_TR COREBCLKSCLKALIGN_0 (.current_state_0(
        current_state_0), .PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE(
        PF_CLK_DIV_FIFO_DELAY_LINE_OUT_OF_RANGE), 
        .PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE(
        PF_IOD_GENERIC_RX_C1_0_CLK_TRAIN_DONE), .CLK_TRAIN_ERROR_c(
        CLK_TRAIN_ERROR_c), .COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE(
        COREBCLKSCLKALIGN_0_BCLKSCLK_ALGN_PAUSE), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_MOV), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_LOAD), 
        .COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS(
        COREBCLKSCLKALIGN_0_ICB_CLK_ALGN_CLR_FLGS), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_LATE_0), 
        .PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0(
        PF_IOD_CLK_TRAINING_EYE_MONITOR_EARLY_0), 
        .RX_CLK_ALIGN_DONE_arst(RX_CLK_ALIGN_DONE_arst), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G));
    
endmodule


module 
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_TRNG_Z1_0(
        
       BIT_ALGN_EYE_IN_c,
       EYE_MONITOR_EARLY_net_0_0,
       EYE_MONITOR_LATE_net_0_0,
       PLL_LOCK_0,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS,
       BIT_ALGN_DONE_0_c,
       BIT_ALGN_START_0_c,
       BIT_ALGN_OOR_0_c,
       BIT_ALGN_ERR_c,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD,
       debouncer_0_DB_OUT,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst
    );
input  [2:0] BIT_ALGN_EYE_IN_c;
input  EYE_MONITOR_EARLY_net_0_0;
input  EYE_MONITOR_LATE_net_0_0;
input  PLL_LOCK_0;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS;
output BIT_ALGN_DONE_0_c;
output BIT_ALGN_START_0_c;
input  BIT_ALGN_OOR_0_c;
output BIT_ALGN_ERR_c;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD;
input  debouncer_0_DB_OUT;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  RX_CLK_ALIGN_DONE_arst;

    wire [9:0] rst_cnt_Z;
    wire [8:0] rst_cnt_s;
    wire [127:0] late_flags_Z;
    wire [127:0] un10_early_flags;
    wire [127:0] late_flags_7_fast_0;
    wire [50:49] late_flags_RNO_0;
    wire [127:0] early_flags_Z;
    wire [127:0] early_flags_7_fast_0;
    wire [50:49] early_flags_RNO_0;
    wire [3:0] restart_edge_reg_Z;
    wire [2:0] restart_reg_Z;
    wire [6:0] tap_cnt_Z;
    wire [2:0] wait_cnt_Z;
    wire [2:0] wait_cnt_4_Z;
    wire [2:0] retrain_reg_Z;
    wire [1:1] cnt_Z;
    wire [1:1] cnt_RNO_0;
    wire [6:0] tapcnt_final_Z;
    wire [6:0] tapcnt_final_13_1_Z;
    wire [6:0] no_early_no_late_val_st1_Z;
    wire [6:0] emflag_cnt_Z;
    wire [6:0] no_early_no_late_val_end2_Z;
    wire [4:0] bitalign_curr_state_Z;
    wire [4:0] bitalign_curr_state_34;
    wire [7:0] noearly_nolate_diff_nxt_8;
    wire [6:0] tapcnt_final_upd_Z;
    wire [1:0] tapcnt_final_upd_8_Z;
    wire [6:3] tapcnt_final_upd_8;
    wire [6:0] early_val_Z;
    wire [6:0] late_val_Z;
    wire [6:0] no_early_no_late_val_st2_Z;
    wire [7:0] early_late_diff_Z;
    wire [7:0] early_late_diff_8;
    wire [7:0] noearly_nolate_diff_start_7;
    wire [6:0] no_early_no_late_val_end1_Z;
    wire [7:0] timeout_cnt_Z;
    wire [7:0] timeout_cnt_s;
    wire [5:0] emflag_cnt_s;
    wire [6:6] emflag_cnt_s_Z;
    wire [9:9] rst_cnt_s_Z;
    wire [6:0] timeout_cnt_cry;
    wire [0:0] timeout_cnt_RNI9ABM_Y_0;
    wire [1:1] timeout_cnt_RNI8UO41_Y_0;
    wire [2:2] timeout_cnt_RNI8J6J1_Y_0;
    wire [3:3] timeout_cnt_RNI99K12_Y_0;
    wire [4:4] timeout_cnt_RNIB02G2_Y_0;
    wire [5:5] timeout_cnt_RNIEOFU2_Y_0;
    wire [7:7] timeout_cnt_RNO_FCO_0;
    wire [7:7] timeout_cnt_RNO_Y_0;
    wire [6:6] timeout_cnt_RNIIHTC3_Y_0;
    wire [0:0] emflag_cnt_cry_cy_S_1;
    wire [0:0] emflag_cnt_cry_cy_Y_1;
    wire [5:0] emflag_cnt_cry_Z;
    wire [5:0] emflag_cnt_cry_Y_1;
    wire [6:6] emflag_cnt_s_FCO_0;
    wire [6:6] emflag_cnt_s_Y_0;
    wire [0:0] un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_S_0;
    wire [0:0] un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_Y_0;
    wire [1:1] tapcnt_final_RNIOTM22_Y_0;
    wire [1:1] un1_tap_cnt_0_sqmuxa_14_0_0;
    wire [2:2] tapcnt_final_RNI2SF33_Y_0;
    wire [3:3] tapcnt_final_RNIES844_Y_0;
    wire [4:4] tapcnt_final_RNISU155_Y_0;
    wire [6:6] tap_cnt_RNO_0_FCO_0;
    wire [6:6] tap_cnt_RNO_0_Y_0;
    wire [5:5] tapcnt_final_RNIC3R56_Y_0;
    wire [0:0] early_val_RNIBEUF3_S;
    wire [0:0] early_val_RNIBEUF3_Y;
    wire [0:0] early_val_RNIT5J81_Z;
    wire [0:0] un1_no_early_no_late_val_end1_1_1_RNIHEIR_0;
    wire [6:1] tapcnt_final_13_m1;
    wire [1:1] early_val_RNIS2TV6_Y;
    wire [1:1] early_val_RNI09J81_Z;
    wire [1:1] un1_no_early_no_late_val_end1_1_1_RNIJGIR_0;
    wire [2:2] early_val_RNIJTRFA_Y;
    wire [2:2] early_val_RNI3CJ81_Z;
    wire [2:2] un1_no_early_no_late_val_end1_1_1_RNILIIR_0;
    wire [3:3] early_val_RNIGUQVD_Y;
    wire [3:3] early_val_RNI6FJ81_Z;
    wire [3:3] un1_no_early_no_late_val_end1_1_1_RNINKIR_0;
    wire [4:4] early_val_RNIJ5QFH_Y;
    wire [4:4] early_val_RNI9IJ81_Z;
    wire [4:4] un1_no_early_no_late_val_end1_1_1_RNIPMIR_0;
    wire [6:6] tapcnt_final_13_RNO_FCO_0;
    wire [6:6] tapcnt_final_13_RNO_Y_0;
    wire [5:5] early_val_RNISIPVK_Y;
    wire [5:5] early_val_RNICLJ81_Z;
    wire [5:5] un1_no_early_no_late_val_end1_1_1_RNIROIR_0;
    wire [8:1] rst_cnt_cry_Z;
    wire [8:1] rst_cnt_cry_Y_1;
    wire [9:9] rst_cnt_s_FCO_1;
    wire [9:9] rst_cnt_s_Y_1;
    wire [6:1] tapcnt_final_13_Z;
    wire [96:0] un10_early_flags_1_Z;
    wire [69:0] un10_early_flags_2_Z;
    wire [100:0] un10_early_flags_2_0;
    wire [87:46] un10_early_flags_3_Z;
    wire [127:127] early_flags_dec;
    wire [6:0] un1_no_early_no_late_val_end1_1_1_Z;
    wire [6:0] un1_no_early_no_late_val_st1_1_1;
    wire [0:0] tapcnt_final_13_1_1_0_Z;
    wire [15:15] un10_early_flags_1_0;
    wire mv_dn_fg_0_sqmuxa_i_o2_0, N_12_i, CO0_0, CO0_0_i, 
        un1_restart_trng_fg_5_0, N_19_i, N_209, N_208, VCC, GND, 
        N_28_i, N_26_i, N_24_i, N_1497_i, N_1496_i, sig_re_train_Z, 
        Restart_trng_edge_det_Z, N_32_i, N_30_i, 
        no_early_no_late_val_st1_0_sqmuxa_i_Z, 
        no_early_no_late_val_end2_0_sqmuxa_i, un16_tapcnt_final_4, 
        un16_tapcnt_final_5, un16_tapcnt_final_6, un16_tapcnt_final_7, 
        tapcnt_final_upd_0_sqmuxa_i_Z, tapcnt_final_upd_8_cry_2_0_Y_0, 
        early_flags_0_sqmuxa_2_i, early_val_0_sqmuxa_1_i_Z, 
        un16_tapcnt_final_0, un16_tapcnt_final_1, un16_tapcnt_final_2, 
        un16_tapcnt_final_3, early_late_diff_0_sqmuxa_1_i, 
        un1_restart_trng_fg_8_0, un10_tapcnt_final_4, 
        no_early_no_late_val_end1_0_sqmuxa_1_i, un10_tapcnt_final_5, 
        un10_tapcnt_final_6, un10_tapcnt_final_7, un10_tapcnt_final_0, 
        un10_tapcnt_final_1, un10_tapcnt_final_2, un10_tapcnt_final_3, 
        bit_align_start_Z, N_1439_i, bit_align_done_0_sqmuxa_3_i_Z, 
        bit_align_done_Z, bit_align_done_2_sqmuxa_Z, calc_done_Z, 
        N_1431_i, calc_done_0_sqmuxa_2_i_Z, rx_trng_done1_Z, N_1415_i, 
        rx_trng_done1_0_sqmuxa_i_Z, rx_BIT_ALGN_LOAD_9, 
        rx_BIT_ALGN_LOAD_0_sqmuxa_1_i_Z, late_last_set_Z, 
        early_late_diff_2_sqmuxa_Z, un1_restart_trng_fg_6_Z, 
        rx_BIT_ALGN_DIR_0_sqmuxa_2_i_Z, rx_BIT_ALGN_MOVE_2_sqmuxa_Z, 
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_i_Z, bit_align_dly_done_Z, 
        bit_align_dly_done_2_sqmuxa_Z, 
        bit_align_dly_done_0_sqmuxa_1_i_Z, rx_trng_done_Z, N_1403, 
        rx_trng_done_0_sqmuxa_i_Z, reset_dly_fg_Z, reset_dly_fg4_Z, 
        sig_rx_BIT_ALGN_CLR_FLGS_Z, sig_rx_BIT_ALGN_CLR_FLGS_11, 
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i_Z, rx_err_Z, N_1392, 
        rx_err_0_sqmuxa_1_i_Z, late_cur_set_Z, late_cur_set_2_sqmuxa, 
        late_cur_set_0_sqmuxa_i, early_cur_set_Z, early_val_2_sqmuxa_Z, 
        early_cur_set_0_sqmuxa_i_Z, early_last_set_Z, 
        early_last_set_2_sqmuxa_Z, early_last_set_0_sqmuxa_i_Z, 
        mv_up_fg_Z, tapcnt_final_upd_2_sqmuxa_1, 
        mv_up_fg_0_sqmuxa_i_0_0, mv_dn_fg_Z, 
        tapcnt_final_upd_3_sqmuxa_1, mv_dn_fg_0_sqmuxa_i_0_0, 
        timeout_cnte, emflag_cnte, timeout_cnt_cry_cy, 
        restart_trng_fg_RNIBNT7_S_0, restart_trng_fg_RNIBNT7_Y_0, 
        restart_trng_fg_i, emflag_cnt_cry_cy, 
        un1_restart_trng_fg_9_0_443_0, 
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Z, 
        noearly_nolate_diff_nxt_8_cry_0_0_cy_S_0, 
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Y_0, 
        noearly_nolate_diff_nxt_8_cry_0, 
        noearly_nolate_diff_nxt_8_cry_0_0_Y_0, 
        noearly_nolate_diff_nxt_8_cry_1, 
        noearly_nolate_diff_nxt_8_cry_1_0_Y_0, 
        noearly_nolate_diff_nxt_8_cry_2, 
        noearly_nolate_diff_nxt_8_cry_2_0_Y_0, 
        noearly_nolate_diff_nxt_8_cry_3, 
        noearly_nolate_diff_nxt_8_cry_3_0_Y_0, 
        noearly_nolate_diff_nxt_8_cry_4, 
        noearly_nolate_diff_nxt_8_cry_4_0_Y_0, 
        noearly_nolate_diff_nxt_8_cry_5, 
        noearly_nolate_diff_nxt_8_cry_5_0_Y_0, 
        noearly_nolate_diff_nxt_8_s_7_FCO_0, 
        noearly_nolate_diff_nxt_8_s_7_Y_0, 
        noearly_nolate_diff_nxt_8_cry_6, 
        noearly_nolate_diff_nxt_8_cry_6_0_Y_0, 
        early_late_diff_8_cry_0_0_cy_Z, 
        early_late_diff_8_cry_0_0_cy_S_0, 
        early_late_diff_8_cry_0_0_cy_Y_0, early_late_diff_8_cry_0, 
        early_late_diff_8_cry_0_0_Y_0, early_late_diff_8_cry_1, 
        early_late_diff_8_cry_1_0_Y_0, early_late_diff_8_cry_2, 
        early_late_diff_8_cry_2_0_Y_0, early_late_diff_8_cry_3, 
        early_late_diff_8_cry_3_0_Y_0, early_late_diff_8_cry_4, 
        early_late_diff_8_cry_4_0_Y_0, early_late_diff_8_cry_5, 
        early_late_diff_8_cry_5_0_Y_0, early_late_diff_8_s_7_FCO_0, 
        early_late_diff_8_s_7_Y_0, early_late_diff_8_cry_6, 
        early_late_diff_8_cry_6_0_Y_0, 
        noearly_nolate_diff_start_7_cry_0_0_cy_Z, 
        noearly_nolate_diff_start_7_cry_0_0_cy_S_0, 
        noearly_nolate_diff_start_7_cry_0_0_cy_Y_0, 
        noearly_nolate_diff_start_7_cry_0, 
        noearly_nolate_diff_start_7_cry_0_0_Y_0, 
        noearly_nolate_diff_start_7_cry_1, 
        noearly_nolate_diff_start_7_cry_1_0_Y_0, 
        noearly_nolate_diff_start_7_cry_2, 
        noearly_nolate_diff_start_7_cry_2_0_Y_0, 
        noearly_nolate_diff_start_7_cry_3, 
        noearly_nolate_diff_start_7_cry_3_0_Y_0, 
        noearly_nolate_diff_start_7_cry_4, 
        noearly_nolate_diff_start_7_cry_4_0_Y_0, 
        noearly_nolate_diff_start_7_cry_5, 
        noearly_nolate_diff_start_7_cry_5_0_Y_0, 
        noearly_nolate_diff_start_7_s_7_FCO_0, 
        noearly_nolate_diff_start_7_s_7_Y_0, 
        noearly_nolate_diff_start_7_cry_6, 
        noearly_nolate_diff_start_7_cry_6_0_Y_0, tap_cnt_17_i_m2_cry_0, 
        N_60, N_89, tap_cnt_17_i_m2_cry_1, N_79, tap_cnt_17_i_m2_cry_2, 
        N_78, tap_cnt_17_i_m2_cry_3, N_77, tap_cnt_17_i_m2_cry_4, N_76, 
        N_74, tap_cnt_17_i_m2_cry_5, N_75, tapcnt_final_13_m1_cry_0, 
        un1_bitalign_curr_state169_12_sn, tapcnt_final_13_m1_cry_1, 
        tapcnt_final_13_m1_cry_2, tapcnt_final_13_m1_cry_3, 
        tapcnt_final_13_m1_cry_4, tapcnt_final_3_sqmuxa_Z, 
        tapcnt_final_13_m1_axb_6_1, tapcnt_final_13_m1_cry_5, 
        tapcnt_final_upd_8_cry_2, tapcnt_final_upd_8_cry_2_0_S_0, 
        tapcnt_final_upd_1_sqmuxa, tapcnt_final_upd_8_cry_3, 
        tapcnt_final_upd_8_cry_3_0_Y_0, tapcnt_final_upd_8_cry_4, 
        tapcnt_final_upd_8_cry_4_0_Y_0, tapcnt_final_upd_8_s_6_FCO_0, 
        tapcnt_final_upd_8_s_6_Y_0, tapcnt_final_upd_8_cry_5, 
        tapcnt_final_upd_8_cry_5_0_Y_0, tapcnt_final27_cry_0_Z, 
        tapcnt_final27_cry_0_S_0, tapcnt_final27_cry_0_Y_0, 
        tapcnt_final27_cry_1_Z, tapcnt_final27_cry_1_S_0, 
        tapcnt_final27_cry_1_Y_0, tapcnt_final27_cry_2_Z, 
        tapcnt_final27_cry_2_S_0, tapcnt_final27_cry_2_Y_0, 
        tapcnt_final27_cry_3_Z, tapcnt_final27_cry_3_S_0, 
        tapcnt_final27_cry_3_Y_0, tapcnt_final27_cry_4_Z, 
        tapcnt_final27_cry_4_S_0, tapcnt_final27_cry_4_Y_0, 
        tapcnt_final27_cry_5_Z, tapcnt_final27_cry_5_S_0, 
        tapcnt_final27_cry_5_Y_0, tapcnt_final27, 
        tapcnt_final27_cry_6_S_0, tapcnt_final27_cry_6_Y_0, 
        un16_tapcnt_final_cry_0_Z, un16_tapcnt_final_cry_0_S_0, 
        un16_tapcnt_final_cry_0_Y_0, un16_tapcnt_final_cry_1_Z, 
        un16_tapcnt_final_cry_1_S_0, un16_tapcnt_final_cry_1_Y_0, 
        un16_tapcnt_final_cry_2_Z, un16_tapcnt_final_cry_2_S_0, 
        un16_tapcnt_final_cry_2_Y_0, un16_tapcnt_final_cry_3_Z, 
        un16_tapcnt_final_cry_3_S_0, un16_tapcnt_final_cry_3_Y_0, 
        un16_tapcnt_final_cry_4_Z, un16_tapcnt_final_cry_4_S_0, 
        un16_tapcnt_final_cry_4_Y_0, un16_tapcnt_final_cry_5_Z, 
        un16_tapcnt_final_cry_5_S_0, un16_tapcnt_final_cry_5_Y_0, 
        un16_tapcnt_final_cry_6_Z, un16_tapcnt_final_cry_6_S_0, 
        un16_tapcnt_final_cry_6_Y_0, un16_tapcnt_final_cry_7_Z, 
        un16_tapcnt_final_cry_7_S_0, un16_tapcnt_final_cry_7_Y_0, 
        un1_early_late_diff_1_cry_0_Z, un1_early_late_diff_1_cry_0_S_0, 
        un1_early_late_diff_1_cry_0_Y_0, un1_early_late_diff_1_cry_1_Z, 
        un1_early_late_diff_1_cry_1_S_0, 
        un1_early_late_diff_1_cry_1_Y_0, un1_early_late_diff_1_cry_2_Z, 
        un1_early_late_diff_1_cry_2_S_0, 
        un1_early_late_diff_1_cry_2_Y_0, un1_early_late_diff_1_cry_3_Z, 
        un1_early_late_diff_1_cry_3_S_0, 
        un1_early_late_diff_1_cry_3_Y_0, un1_early_late_diff_1_cry_4_Z, 
        un1_early_late_diff_1_cry_4_S_0, 
        un1_early_late_diff_1_cry_4_Y_0, un1_early_late_diff_1_cry_5_Z, 
        un1_early_late_diff_1_cry_5_S_0, 
        un1_early_late_diff_1_cry_5_Y_0, un1_early_late_diff_1_cry_6_Z, 
        un1_early_late_diff_1_cry_6_S_0, 
        un1_early_late_diff_1_cry_6_Y_0, un1_early_late_diff_1_cry_7_Z, 
        un1_early_late_diff_1_cry_7_S_0, 
        un1_early_late_diff_1_cry_7_Y_0, un10_tapcnt_final_cry_0_Z, 
        un10_tapcnt_final_cry_0_S_0, un10_tapcnt_final_cry_0_Y_0, 
        un10_tapcnt_final_cry_1_Z, un10_tapcnt_final_cry_1_S_0, 
        un10_tapcnt_final_cry_1_Y_0, un10_tapcnt_final_cry_2_Z, 
        un10_tapcnt_final_cry_2_S_0, un10_tapcnt_final_cry_2_Y_0, 
        un10_tapcnt_final_cry_3_Z, un10_tapcnt_final_cry_3_S_0, 
        un10_tapcnt_final_cry_3_Y_0, un10_tapcnt_final_cry_4_Z, 
        un10_tapcnt_final_cry_4_S_0, un10_tapcnt_final_cry_4_Y_0, 
        un10_tapcnt_final_cry_5_Z, un10_tapcnt_final_cry_5_S_0, 
        un10_tapcnt_final_cry_5_Y_0, un10_tapcnt_final_cry_6_Z, 
        un10_tapcnt_final_cry_6_S_0, un10_tapcnt_final_cry_6_Y_0, 
        un10_tapcnt_final_cry_7_Z, un10_tapcnt_final_cry_7_S_0, 
        un10_tapcnt_final_cry_7_Y_0, un1_early_late_diff_cry_0_Z, 
        un1_early_late_diff_cry_0_S_0, un1_early_late_diff_cry_0_Y_0, 
        un1_early_late_diff_cry_1_Z, un1_early_late_diff_cry_1_S_0, 
        un1_early_late_diff_cry_1_Y_0, un1_early_late_diff_cry_2_Z, 
        un1_early_late_diff_cry_2_S_0, un1_early_late_diff_cry_2_Y_0, 
        un1_early_late_diff_cry_3_Z, un1_early_late_diff_cry_3_S_0, 
        un1_early_late_diff_cry_3_Y_0, un1_early_late_diff_cry_4_Z, 
        un1_early_late_diff_cry_4_S_0, un1_early_late_diff_cry_4_Y_0, 
        un1_early_late_diff_cry_5_Z, un1_early_late_diff_cry_5_S_0, 
        un1_early_late_diff_cry_5_Y_0, un1_early_late_diff_cry_6_Z, 
        un1_early_late_diff_cry_6_S_0, un1_early_late_diff_cry_6_Y_0, 
        un1_early_late_diff_cry_7_Z, un1_early_late_diff_cry_7_S_0, 
        un1_early_late_diff_cry_7_Y_0, rst_cnt_s_715_FCO_0, 
        rst_cnt_s_715_S_0, rst_cnt_s_715_Y_0, 
        late_flags_pmux_127_1_0_co1, 
        late_flags_pmux_127_1_0_wmux_0_S_0, late_flags_pmux, 
        late_flags_pmux_126_1_1_wmux_10_Y_0, 
        late_flags_pmux_126_1_0_wmux_10_Y_0, 
        late_flags_pmux_127_1_0_y0, late_flags_pmux_127_1_0_co0, 
        late_flags_pmux_127_1_0_wmux_S_0, 
        late_flags_pmux_63_1_1_wmux_10_Y_0, 
        late_flags_pmux_63_1_0_wmux_10_Y_0, 
        early_flags_pmux_127_1_0_co1, 
        early_flags_pmux_127_1_0_wmux_0_S_0, early_flags_pmux, 
        early_flags_pmux_126_1_1_wmux_10_Y_0, 
        early_flags_pmux_126_1_0_wmux_10_Y_0, 
        early_flags_pmux_127_1_0_y0, early_flags_pmux_127_1_0_co0, 
        early_flags_pmux_127_1_0_wmux_S_0, 
        early_flags_pmux_63_1_1_wmux_10_Y_0, 
        early_flags_pmux_63_1_0_wmux_10_Y_0, m74_2_1_1_1_co1, 
        m74_2_1_1_wmux_0_S_0, N_75_0, N_29_i, N_116_mux, 
        m74_2_1_1_1_y0, m74_2_1_1_1_co0, m74_2_1_1_wmux_S_0, N_69, 
        m74_1_0_0, early_flags_pmux_63_1_1_co1_9, 
        early_flags_pmux_63_1_1_wmux_20_S_0, 
        early_flags_pmux_63_1_1_y21, early_flags_pmux_63_1_1_y3_0, 
        early_flags_pmux_63_1_1_y1_0, early_flags_pmux_63_1_1_y0_8, 
        early_flags_pmux_63_1_1_co0_9, 
        early_flags_pmux_63_1_1_wmux_19_S_0, 
        early_flags_pmux_63_1_1_y5_0, early_flags_pmux_63_1_1_y7_0, 
        early_flags_pmux_63_1_1_co1_8, 
        early_flags_pmux_63_1_1_wmux_18_S_0, 
        early_flags_pmux_63_1_1_y0_7, early_flags_pmux_63_1_1_co0_8, 
        early_flags_pmux_63_1_1_wmux_17_S_0, 
        early_flags_pmux_63_1_1_co1_7, 
        early_flags_pmux_63_1_1_wmux_16_S_0, 
        early_flags_pmux_63_1_1_y0_6, early_flags_pmux_63_1_1_co0_7, 
        early_flags_pmux_63_1_1_wmux_15_S_0, 
        early_flags_pmux_63_1_1_co1_6, 
        early_flags_pmux_63_1_1_wmux_14_S_0, 
        early_flags_pmux_63_1_1_y0_5, early_flags_pmux_63_1_1_co0_6, 
        early_flags_pmux_63_1_1_wmux_13_S_0, 
        early_flags_pmux_63_1_1_co1_5, 
        early_flags_pmux_63_1_1_wmux_12_S_0, 
        early_flags_pmux_63_1_1_y0_4, early_flags_pmux_63_1_1_co0_5, 
        early_flags_pmux_63_1_1_wmux_11_S_0, 
        early_flags_pmux_63_1_1_co1_4, 
        early_flags_pmux_63_1_1_wmux_10_S_0, 
        early_flags_pmux_63_1_1_y9, early_flags_pmux_63_1_1_co0_4, 
        early_flags_pmux_63_1_1_wmux_9_S_0, 
        early_flags_pmux_63_1_1_wmux_9_Y_0, 
        early_flags_pmux_63_1_1_co1_3, 
        early_flags_pmux_63_1_1_wmux_8_S_0, early_flags_pmux_63_1_1_y3, 
        early_flags_pmux_63_1_1_y1, early_flags_pmux_63_1_1_y0_3, 
        early_flags_pmux_63_1_1_co0_3, 
        early_flags_pmux_63_1_1_wmux_7_S_0, early_flags_pmux_63_1_1_y5, 
        early_flags_pmux_63_1_1_y7, early_flags_pmux_63_1_1_co1_2, 
        early_flags_pmux_63_1_1_wmux_6_S_0, 
        early_flags_pmux_63_1_1_y0_2, early_flags_pmux_63_1_1_co0_2, 
        early_flags_pmux_63_1_1_wmux_5_S_0, 
        early_flags_pmux_63_1_1_co1_1, 
        early_flags_pmux_63_1_1_wmux_4_S_0, 
        early_flags_pmux_63_1_1_y0_1, early_flags_pmux_63_1_1_co0_1, 
        early_flags_pmux_63_1_1_wmux_3_S_0, 
        early_flags_pmux_63_1_1_co1_0, 
        early_flags_pmux_63_1_1_wmux_2_S_0, 
        early_flags_pmux_63_1_1_y0_0, early_flags_pmux_63_1_1_co0_0, 
        early_flags_pmux_63_1_1_wmux_1_S_0, 
        early_flags_pmux_63_1_1_co1, 
        early_flags_pmux_63_1_1_wmux_0_S_0, early_flags_pmux_63_1_1_y0, 
        early_flags_pmux_63_1_1_co0, early_flags_pmux_63_1_1_wmux_S_0, 
        late_flags_pmux_126_1_1_co1_9, 
        late_flags_pmux_126_1_1_wmux_20_S_0, 
        late_flags_pmux_126_1_1_y21, late_flags_pmux_126_1_1_y3_0, 
        late_flags_pmux_126_1_1_y1_0, late_flags_pmux_126_1_1_y0_8, 
        late_flags_pmux_126_1_1_co0_9, 
        late_flags_pmux_126_1_1_wmux_19_S_0, 
        late_flags_pmux_126_1_1_y5_0, late_flags_pmux_126_1_1_y7_0, 
        late_flags_pmux_126_1_1_co1_8, 
        late_flags_pmux_126_1_1_wmux_18_S_0, 
        late_flags_pmux_126_1_1_y0_7, late_flags_pmux_126_1_1_co0_8, 
        late_flags_pmux_126_1_1_wmux_17_S_0, 
        late_flags_pmux_126_1_1_co1_7, 
        late_flags_pmux_126_1_1_wmux_16_S_0, 
        late_flags_pmux_126_1_1_y0_6, late_flags_pmux_126_1_1_co0_7, 
        late_flags_pmux_126_1_1_wmux_15_S_0, 
        late_flags_pmux_126_1_1_co1_6, 
        late_flags_pmux_126_1_1_wmux_14_S_0, 
        late_flags_pmux_126_1_1_y0_5, late_flags_pmux_126_1_1_co0_6, 
        late_flags_pmux_126_1_1_wmux_13_S_0, 
        late_flags_pmux_126_1_1_co1_5, 
        late_flags_pmux_126_1_1_wmux_12_S_0, 
        late_flags_pmux_126_1_1_y0_4, late_flags_pmux_126_1_1_co0_5, 
        late_flags_pmux_126_1_1_wmux_11_S_0, 
        late_flags_pmux_126_1_1_co1_4, 
        late_flags_pmux_126_1_1_wmux_10_S_0, 
        late_flags_pmux_126_1_1_y9, late_flags_pmux_126_1_1_co0_4, 
        late_flags_pmux_126_1_1_wmux_9_S_0, 
        late_flags_pmux_126_1_1_wmux_9_Y_0, 
        late_flags_pmux_126_1_1_co1_3, 
        late_flags_pmux_126_1_1_wmux_8_S_0, late_flags_pmux_126_1_1_y3, 
        late_flags_pmux_126_1_1_y1, late_flags_pmux_126_1_1_y0_3, 
        late_flags_pmux_126_1_1_co0_3, 
        late_flags_pmux_126_1_1_wmux_7_S_0, late_flags_pmux_126_1_1_y5, 
        late_flags_pmux_126_1_1_y7, late_flags_pmux_126_1_1_co1_2, 
        late_flags_pmux_126_1_1_wmux_6_S_0, 
        late_flags_pmux_126_1_1_y0_2, late_flags_pmux_126_1_1_co0_2, 
        late_flags_pmux_126_1_1_wmux_5_S_0, 
        late_flags_pmux_126_1_1_co1_1, 
        late_flags_pmux_126_1_1_wmux_4_S_0, 
        late_flags_pmux_126_1_1_y0_1, late_flags_pmux_126_1_1_co0_1, 
        late_flags_pmux_126_1_1_wmux_3_S_0, 
        late_flags_pmux_126_1_1_co1_0, 
        late_flags_pmux_126_1_1_wmux_2_S_0, 
        late_flags_pmux_126_1_1_y0_0, late_flags_pmux_126_1_1_co0_0, 
        late_flags_pmux_126_1_1_wmux_1_S_0, 
        late_flags_pmux_126_1_1_co1, 
        late_flags_pmux_126_1_1_wmux_0_S_0, late_flags_pmux_126_1_1_y0, 
        late_flags_pmux_126_1_1_co0, late_flags_pmux_126_1_1_wmux_S_0, 
        late_flags_pmux_63_1_0_co1_9, 
        late_flags_pmux_63_1_0_wmux_20_S_0, 
        late_flags_pmux_63_1_0_0_y21, late_flags_pmux_63_1_0_y3_0, 
        late_flags_pmux_63_1_0_y1_0, late_flags_pmux_63_1_0_y0_8, 
        late_flags_pmux_63_1_0_co0_9, 
        late_flags_pmux_63_1_0_wmux_19_S_0, 
        late_flags_pmux_63_1_0_y5_0, late_flags_pmux_63_1_0_y7_0, 
        late_flags_pmux_63_1_0_co1_8, 
        late_flags_pmux_63_1_0_wmux_18_S_0, 
        late_flags_pmux_63_1_0_y0_7, late_flags_pmux_63_1_0_co0_8, 
        late_flags_pmux_63_1_0_wmux_17_S_0, 
        late_flags_pmux_63_1_0_co1_7, 
        late_flags_pmux_63_1_0_wmux_16_S_0, 
        late_flags_pmux_63_1_0_y0_6, late_flags_pmux_63_1_0_co0_7, 
        late_flags_pmux_63_1_0_wmux_15_S_0, 
        late_flags_pmux_63_1_0_co1_6, 
        late_flags_pmux_63_1_0_wmux_14_S_0, 
        late_flags_pmux_63_1_0_y0_5, late_flags_pmux_63_1_0_co0_6, 
        late_flags_pmux_63_1_0_wmux_13_S_0, 
        late_flags_pmux_63_1_0_co1_5, 
        late_flags_pmux_63_1_0_wmux_12_S_0, 
        late_flags_pmux_63_1_0_y0_4, late_flags_pmux_63_1_0_co0_5, 
        late_flags_pmux_63_1_0_wmux_11_S_0, 
        late_flags_pmux_63_1_0_co1_4, 
        late_flags_pmux_63_1_0_wmux_10_S_0, 
        late_flags_pmux_63_1_0_0_y9, late_flags_pmux_63_1_0_co0_4, 
        late_flags_pmux_63_1_0_wmux_9_S_0, 
        late_flags_pmux_63_1_0_wmux_9_Y_0, 
        late_flags_pmux_63_1_0_co1_3, 
        late_flags_pmux_63_1_0_wmux_8_S_0, late_flags_pmux_63_1_0_0_y3, 
        late_flags_pmux_63_1_0_0_y1, late_flags_pmux_63_1_0_y0_3, 
        late_flags_pmux_63_1_0_co0_3, 
        late_flags_pmux_63_1_0_wmux_7_S_0, late_flags_pmux_63_1_0_0_y5, 
        late_flags_pmux_63_1_0_0_y7, late_flags_pmux_63_1_0_co1_2, 
        late_flags_pmux_63_1_0_wmux_6_S_0, late_flags_pmux_63_1_0_y0_2, 
        late_flags_pmux_63_1_0_co0_2, 
        late_flags_pmux_63_1_0_wmux_5_S_0, 
        late_flags_pmux_63_1_0_co1_1, 
        late_flags_pmux_63_1_0_wmux_4_S_0, late_flags_pmux_63_1_0_y0_1, 
        late_flags_pmux_63_1_0_co0_1, 
        late_flags_pmux_63_1_0_wmux_3_S_0, 
        late_flags_pmux_63_1_0_co1_0, 
        late_flags_pmux_63_1_0_wmux_2_S_0, late_flags_pmux_63_1_0_y0_0, 
        late_flags_pmux_63_1_0_co0_0, 
        late_flags_pmux_63_1_0_wmux_1_S_0, 
        late_flags_pmux_63_1_0_0_co1, 
        late_flags_pmux_63_1_0_wmux_0_S_0, late_flags_pmux_63_1_0_0_y0, 
        late_flags_pmux_63_1_0_0_co0, late_flags_pmux_63_1_0_wmux_S_0, 
        early_flags_pmux_126_1_0_co1_9, 
        early_flags_pmux_126_1_0_wmux_20_S_0, 
        early_flags_pmux_126_1_0_0_y21, early_flags_pmux_126_1_0_y3_0, 
        early_flags_pmux_126_1_0_y1_0, early_flags_pmux_126_1_0_y0_8, 
        early_flags_pmux_126_1_0_co0_9, 
        early_flags_pmux_126_1_0_wmux_19_S_0, 
        early_flags_pmux_126_1_0_y5_0, early_flags_pmux_126_1_0_y7_0, 
        early_flags_pmux_126_1_0_co1_8, 
        early_flags_pmux_126_1_0_wmux_18_S_0, 
        early_flags_pmux_126_1_0_y0_7, early_flags_pmux_126_1_0_co0_8, 
        early_flags_pmux_126_1_0_wmux_17_S_0, 
        early_flags_pmux_126_1_0_co1_7, 
        early_flags_pmux_126_1_0_wmux_16_S_0, 
        early_flags_pmux_126_1_0_y0_6, early_flags_pmux_126_1_0_co0_7, 
        early_flags_pmux_126_1_0_wmux_15_S_0, 
        early_flags_pmux_126_1_0_co1_6, 
        early_flags_pmux_126_1_0_wmux_14_S_0, 
        early_flags_pmux_126_1_0_y0_5, early_flags_pmux_126_1_0_co0_6, 
        early_flags_pmux_126_1_0_wmux_13_S_0, 
        early_flags_pmux_126_1_0_co1_5, 
        early_flags_pmux_126_1_0_wmux_12_S_0, 
        early_flags_pmux_126_1_0_y0_4, early_flags_pmux_126_1_0_co0_5, 
        early_flags_pmux_126_1_0_wmux_11_S_0, 
        early_flags_pmux_126_1_0_co1_4, 
        early_flags_pmux_126_1_0_wmux_10_S_0, 
        early_flags_pmux_126_1_0_0_y9, early_flags_pmux_126_1_0_co0_4, 
        early_flags_pmux_126_1_0_wmux_9_S_0, 
        early_flags_pmux_126_1_0_wmux_9_Y_0, 
        early_flags_pmux_126_1_0_co1_3, 
        early_flags_pmux_126_1_0_wmux_8_S_0, 
        early_flags_pmux_126_1_0_0_y3, early_flags_pmux_126_1_0_0_y1, 
        early_flags_pmux_126_1_0_y0_3, early_flags_pmux_126_1_0_co0_3, 
        early_flags_pmux_126_1_0_wmux_7_S_0, 
        early_flags_pmux_126_1_0_0_y5, early_flags_pmux_126_1_0_0_y7, 
        early_flags_pmux_126_1_0_co1_2, 
        early_flags_pmux_126_1_0_wmux_6_S_0, 
        early_flags_pmux_126_1_0_y0_2, early_flags_pmux_126_1_0_co0_2, 
        early_flags_pmux_126_1_0_wmux_5_S_0, 
        early_flags_pmux_126_1_0_co1_1, 
        early_flags_pmux_126_1_0_wmux_4_S_0, 
        early_flags_pmux_126_1_0_y0_1, early_flags_pmux_126_1_0_co0_1, 
        early_flags_pmux_126_1_0_wmux_3_S_0, 
        early_flags_pmux_126_1_0_co1_0, 
        early_flags_pmux_126_1_0_wmux_2_S_0, 
        early_flags_pmux_126_1_0_y0_0, early_flags_pmux_126_1_0_co0_0, 
        early_flags_pmux_126_1_0_wmux_1_S_0, 
        early_flags_pmux_126_1_0_0_co1, 
        early_flags_pmux_126_1_0_wmux_0_S_0, 
        early_flags_pmux_126_1_0_0_y0, early_flags_pmux_126_1_0_0_co0, 
        early_flags_pmux_126_1_0_wmux_S_0, 
        early_flags_pmux_126_1_1_co1_9, 
        early_flags_pmux_126_1_1_wmux_20_S_0, 
        early_flags_pmux_126_1_1_y21, early_flags_pmux_126_1_1_y3_0, 
        early_flags_pmux_126_1_1_y1_0, early_flags_pmux_126_1_1_y0_8, 
        early_flags_pmux_126_1_1_co0_9, 
        early_flags_pmux_126_1_1_wmux_19_S_0, 
        early_flags_pmux_126_1_1_y5_0, early_flags_pmux_126_1_1_y7_0, 
        early_flags_pmux_126_1_1_co1_8, 
        early_flags_pmux_126_1_1_wmux_18_S_0, 
        early_flags_pmux_126_1_1_y0_7, early_flags_pmux_126_1_1_co0_8, 
        early_flags_pmux_126_1_1_wmux_17_S_0, 
        early_flags_pmux_126_1_1_co1_7, 
        early_flags_pmux_126_1_1_wmux_16_S_0, 
        early_flags_pmux_126_1_1_y0_6, early_flags_pmux_126_1_1_co0_7, 
        early_flags_pmux_126_1_1_wmux_15_S_0, 
        early_flags_pmux_126_1_1_co1_6, 
        early_flags_pmux_126_1_1_wmux_14_S_0, 
        early_flags_pmux_126_1_1_y0_5, early_flags_pmux_126_1_1_co0_6, 
        early_flags_pmux_126_1_1_wmux_13_S_0, 
        early_flags_pmux_126_1_1_co1_5, 
        early_flags_pmux_126_1_1_wmux_12_S_0, 
        early_flags_pmux_126_1_1_y0_4, early_flags_pmux_126_1_1_co0_5, 
        early_flags_pmux_126_1_1_wmux_11_S_0, 
        early_flags_pmux_126_1_1_co1_4, 
        early_flags_pmux_126_1_1_wmux_10_S_0, 
        early_flags_pmux_126_1_1_y9, early_flags_pmux_126_1_1_co0_4, 
        early_flags_pmux_126_1_1_wmux_9_S_0, 
        early_flags_pmux_126_1_1_wmux_9_Y_0, 
        early_flags_pmux_126_1_1_co1_3, 
        early_flags_pmux_126_1_1_wmux_8_S_0, 
        early_flags_pmux_126_1_1_y3, early_flags_pmux_126_1_1_y1, 
        early_flags_pmux_126_1_1_y0_3, early_flags_pmux_126_1_1_co0_3, 
        early_flags_pmux_126_1_1_wmux_7_S_0, 
        early_flags_pmux_126_1_1_y5, early_flags_pmux_126_1_1_y7, 
        early_flags_pmux_126_1_1_co1_2, 
        early_flags_pmux_126_1_1_wmux_6_S_0, 
        early_flags_pmux_126_1_1_y0_2, early_flags_pmux_126_1_1_co0_2, 
        early_flags_pmux_126_1_1_wmux_5_S_0, 
        early_flags_pmux_126_1_1_co1_1, 
        early_flags_pmux_126_1_1_wmux_4_S_0, 
        early_flags_pmux_126_1_1_y0_1, early_flags_pmux_126_1_1_co0_1, 
        early_flags_pmux_126_1_1_wmux_3_S_0, 
        early_flags_pmux_126_1_1_co1_0, 
        early_flags_pmux_126_1_1_wmux_2_S_0, 
        early_flags_pmux_126_1_1_y0_0, early_flags_pmux_126_1_1_co0_0, 
        early_flags_pmux_126_1_1_wmux_1_S_0, 
        early_flags_pmux_126_1_1_co1, 
        early_flags_pmux_126_1_1_wmux_0_S_0, 
        early_flags_pmux_126_1_1_y0, early_flags_pmux_126_1_1_co0, 
        early_flags_pmux_126_1_1_wmux_S_0, 
        early_flags_pmux_63_1_0_co1_9, 
        early_flags_pmux_63_1_0_wmux_20_S_0, 
        early_flags_pmux_63_1_0_0_y21, early_flags_pmux_63_1_0_y3_0, 
        early_flags_pmux_63_1_0_y1_0, early_flags_pmux_63_1_0_y0_8, 
        early_flags_pmux_63_1_0_co0_9, 
        early_flags_pmux_63_1_0_wmux_19_S_0, 
        early_flags_pmux_63_1_0_y5_0, early_flags_pmux_63_1_0_y7_0, 
        early_flags_pmux_63_1_0_co1_8, 
        early_flags_pmux_63_1_0_wmux_18_S_0, 
        early_flags_pmux_63_1_0_y0_7, early_flags_pmux_63_1_0_co0_8, 
        early_flags_pmux_63_1_0_wmux_17_S_0, 
        early_flags_pmux_63_1_0_co1_7, 
        early_flags_pmux_63_1_0_wmux_16_S_0, 
        early_flags_pmux_63_1_0_y0_6, early_flags_pmux_63_1_0_co0_7, 
        early_flags_pmux_63_1_0_wmux_15_S_0, 
        early_flags_pmux_63_1_0_co1_6, 
        early_flags_pmux_63_1_0_wmux_14_S_0, 
        early_flags_pmux_63_1_0_y0_5, early_flags_pmux_63_1_0_co0_6, 
        early_flags_pmux_63_1_0_wmux_13_S_0, 
        early_flags_pmux_63_1_0_co1_5, 
        early_flags_pmux_63_1_0_wmux_12_S_0, 
        early_flags_pmux_63_1_0_y0_4, early_flags_pmux_63_1_0_co0_5, 
        early_flags_pmux_63_1_0_wmux_11_S_0, 
        early_flags_pmux_63_1_0_co1_4, 
        early_flags_pmux_63_1_0_wmux_10_S_0, 
        early_flags_pmux_63_1_0_0_y9, early_flags_pmux_63_1_0_co0_4, 
        early_flags_pmux_63_1_0_wmux_9_S_0, 
        early_flags_pmux_63_1_0_wmux_9_Y_0, 
        early_flags_pmux_63_1_0_co1_3, 
        early_flags_pmux_63_1_0_wmux_8_S_0, 
        early_flags_pmux_63_1_0_0_y3, early_flags_pmux_63_1_0_0_y1, 
        early_flags_pmux_63_1_0_y0_3, early_flags_pmux_63_1_0_co0_3, 
        early_flags_pmux_63_1_0_wmux_7_S_0, 
        early_flags_pmux_63_1_0_0_y5, early_flags_pmux_63_1_0_0_y7, 
        early_flags_pmux_63_1_0_co1_2, 
        early_flags_pmux_63_1_0_wmux_6_S_0, 
        early_flags_pmux_63_1_0_y0_2, early_flags_pmux_63_1_0_co0_2, 
        early_flags_pmux_63_1_0_wmux_5_S_0, 
        early_flags_pmux_63_1_0_co1_1, 
        early_flags_pmux_63_1_0_wmux_4_S_0, 
        early_flags_pmux_63_1_0_y0_1, early_flags_pmux_63_1_0_co0_1, 
        early_flags_pmux_63_1_0_wmux_3_S_0, 
        early_flags_pmux_63_1_0_co1_0, 
        early_flags_pmux_63_1_0_wmux_2_S_0, 
        early_flags_pmux_63_1_0_y0_0, early_flags_pmux_63_1_0_co0_0, 
        early_flags_pmux_63_1_0_wmux_1_S_0, 
        early_flags_pmux_63_1_0_0_co1, 
        early_flags_pmux_63_1_0_wmux_0_S_0, 
        early_flags_pmux_63_1_0_0_y0, early_flags_pmux_63_1_0_0_co0, 
        early_flags_pmux_63_1_0_wmux_S_0, late_flags_pmux_63_1_1_co1_9, 
        late_flags_pmux_63_1_1_wmux_20_S_0, late_flags_pmux_63_1_1_y21, 
        late_flags_pmux_63_1_1_y3_0, late_flags_pmux_63_1_1_y1_0, 
        late_flags_pmux_63_1_1_y0_8, late_flags_pmux_63_1_1_co0_9, 
        late_flags_pmux_63_1_1_wmux_19_S_0, 
        late_flags_pmux_63_1_1_y5_0, late_flags_pmux_63_1_1_y7_0, 
        late_flags_pmux_63_1_1_co1_8, 
        late_flags_pmux_63_1_1_wmux_18_S_0, 
        late_flags_pmux_63_1_1_y0_7, late_flags_pmux_63_1_1_co0_8, 
        late_flags_pmux_63_1_1_wmux_17_S_0, 
        late_flags_pmux_63_1_1_co1_7, 
        late_flags_pmux_63_1_1_wmux_16_S_0, 
        late_flags_pmux_63_1_1_y0_6, late_flags_pmux_63_1_1_co0_7, 
        late_flags_pmux_63_1_1_wmux_15_S_0, 
        late_flags_pmux_63_1_1_co1_6, 
        late_flags_pmux_63_1_1_wmux_14_S_0, 
        late_flags_pmux_63_1_1_y0_5, late_flags_pmux_63_1_1_co0_6, 
        late_flags_pmux_63_1_1_wmux_13_S_0, 
        late_flags_pmux_63_1_1_co1_5, 
        late_flags_pmux_63_1_1_wmux_12_S_0, 
        late_flags_pmux_63_1_1_y0_4, late_flags_pmux_63_1_1_co0_5, 
        late_flags_pmux_63_1_1_wmux_11_S_0, 
        late_flags_pmux_63_1_1_co1_4, 
        late_flags_pmux_63_1_1_wmux_10_S_0, late_flags_pmux_63_1_1_y9, 
        late_flags_pmux_63_1_1_co0_4, 
        late_flags_pmux_63_1_1_wmux_9_S_0, 
        late_flags_pmux_63_1_1_wmux_9_Y_0, 
        late_flags_pmux_63_1_1_co1_3, 
        late_flags_pmux_63_1_1_wmux_8_S_0, late_flags_pmux_63_1_1_y3, 
        late_flags_pmux_63_1_1_y1, late_flags_pmux_63_1_1_y0_3, 
        late_flags_pmux_63_1_1_co0_3, 
        late_flags_pmux_63_1_1_wmux_7_S_0, late_flags_pmux_63_1_1_y5, 
        late_flags_pmux_63_1_1_y7, late_flags_pmux_63_1_1_co1_2, 
        late_flags_pmux_63_1_1_wmux_6_S_0, late_flags_pmux_63_1_1_y0_2, 
        late_flags_pmux_63_1_1_co0_2, 
        late_flags_pmux_63_1_1_wmux_5_S_0, 
        late_flags_pmux_63_1_1_co1_1, 
        late_flags_pmux_63_1_1_wmux_4_S_0, late_flags_pmux_63_1_1_y0_1, 
        late_flags_pmux_63_1_1_co0_1, 
        late_flags_pmux_63_1_1_wmux_3_S_0, 
        late_flags_pmux_63_1_1_co1_0, 
        late_flags_pmux_63_1_1_wmux_2_S_0, late_flags_pmux_63_1_1_y0_0, 
        late_flags_pmux_63_1_1_co0_0, 
        late_flags_pmux_63_1_1_wmux_1_S_0, late_flags_pmux_63_1_1_co1, 
        late_flags_pmux_63_1_1_wmux_0_S_0, late_flags_pmux_63_1_1_y0, 
        late_flags_pmux_63_1_1_co0, late_flags_pmux_63_1_1_wmux_S_0, 
        late_flags_pmux_126_1_0_co1_9, 
        late_flags_pmux_126_1_0_wmux_20_S_0, 
        late_flags_pmux_126_1_0_0_y21, late_flags_pmux_126_1_0_y3_0, 
        late_flags_pmux_126_1_0_y1_0, late_flags_pmux_126_1_0_y0_8, 
        late_flags_pmux_126_1_0_co0_9, 
        late_flags_pmux_126_1_0_wmux_19_S_0, 
        late_flags_pmux_126_1_0_y5_0, late_flags_pmux_126_1_0_y7_0, 
        late_flags_pmux_126_1_0_co1_8, 
        late_flags_pmux_126_1_0_wmux_18_S_0, 
        late_flags_pmux_126_1_0_y0_7, late_flags_pmux_126_1_0_co0_8, 
        late_flags_pmux_126_1_0_wmux_17_S_0, 
        late_flags_pmux_126_1_0_co1_7, 
        late_flags_pmux_126_1_0_wmux_16_S_0, 
        late_flags_pmux_126_1_0_y0_6, late_flags_pmux_126_1_0_co0_7, 
        late_flags_pmux_126_1_0_wmux_15_S_0, 
        late_flags_pmux_126_1_0_co1_6, 
        late_flags_pmux_126_1_0_wmux_14_S_0, 
        late_flags_pmux_126_1_0_y0_5, late_flags_pmux_126_1_0_co0_6, 
        late_flags_pmux_126_1_0_wmux_13_S_0, 
        late_flags_pmux_126_1_0_co1_5, 
        late_flags_pmux_126_1_0_wmux_12_S_0, 
        late_flags_pmux_126_1_0_y0_4, late_flags_pmux_126_1_0_co0_5, 
        late_flags_pmux_126_1_0_wmux_11_S_0, 
        late_flags_pmux_126_1_0_co1_4, 
        late_flags_pmux_126_1_0_wmux_10_S_0, 
        late_flags_pmux_126_1_0_0_y9, late_flags_pmux_126_1_0_co0_4, 
        late_flags_pmux_126_1_0_wmux_9_S_0, 
        late_flags_pmux_126_1_0_wmux_9_Y_0, 
        late_flags_pmux_126_1_0_co1_3, 
        late_flags_pmux_126_1_0_wmux_8_S_0, 
        late_flags_pmux_126_1_0_0_y3, late_flags_pmux_126_1_0_0_y1, 
        late_flags_pmux_126_1_0_y0_3, late_flags_pmux_126_1_0_co0_3, 
        late_flags_pmux_126_1_0_wmux_7_S_0, 
        late_flags_pmux_126_1_0_0_y5, late_flags_pmux_126_1_0_0_y7, 
        late_flags_pmux_126_1_0_co1_2, 
        late_flags_pmux_126_1_0_wmux_6_S_0, 
        late_flags_pmux_126_1_0_y0_2, late_flags_pmux_126_1_0_co0_2, 
        late_flags_pmux_126_1_0_wmux_5_S_0, 
        late_flags_pmux_126_1_0_co1_1, 
        late_flags_pmux_126_1_0_wmux_4_S_0, 
        late_flags_pmux_126_1_0_y0_1, late_flags_pmux_126_1_0_co0_1, 
        late_flags_pmux_126_1_0_wmux_3_S_0, 
        late_flags_pmux_126_1_0_co1_0, 
        late_flags_pmux_126_1_0_wmux_2_S_0, 
        late_flags_pmux_126_1_0_y0_0, late_flags_pmux_126_1_0_co0_0, 
        late_flags_pmux_126_1_0_wmux_1_S_0, 
        late_flags_pmux_126_1_0_0_co1, 
        late_flags_pmux_126_1_0_wmux_0_S_0, 
        late_flags_pmux_126_1_0_0_y0, late_flags_pmux_126_1_0_0_co0, 
        late_flags_pmux_126_1_0_wmux_S_0, un1_bitalign_curr_state_12_Z, 
        un1_restart_trng_fg_10_sn, un1_retrain_adj_tap_i, 
        un1_rx_BIT_ALGN_START, bitalign_curr_state148_Z, 
        bitalign_curr_state12_Z, bitalign_curr_state_0_sqmuxa_10, 
        bitalign_curr_state160_Z, emflag_cnt_0_sqmuxa, 
        bitalign_curr_state159, un1_early_last_set_1_sqmuxa_1_1_tz_Z, 
        bitalign_curr_state149_Z, tap_cnt_0_sqmuxa_1_Z, 
        sig_rx_BIT_ALGN_CLR_FLGS14_Z, un1_tap_cnt_0_sqmuxa_6_0, 
        un2_noearly_nolate_diff_start_valid, calc_done25, 
        un1_tapcnt_final, calc_done27, bitalign_curr_state162_Z, 
        un1_calc_done25_5, un1_early_late_diff_valid_Z, 
        un10_early_flags_47_0_Z, un10_early_flags_30_0_Z, N_20, 
        late_last_set15_Z, N_94, N_60_0, bitalign_curr_state148_2_Z, 
        N_40, m40_1_1, un1_restart_trng_fg_10_sn_1, 
        early_last_set_1_sqmuxa_1_3_Z, early_val_0_sqmuxa_1_0_Z, N_100, 
        m101_1_1, N_102, bitalign_curr_state161_2_Z, N_92, 
        calc_done25_236, calc_done25_237, calc_done25_253_1_0, 
        calc_done25_245, calc_done25_253, calc_done25_239, 
        calc_done25_238, calc_done25_233, calc_done25_232, m91_1, 
        m91_1_0, m64_1_1, N_63, N_65, bitalign_curr_state41_Z, m82_1_0, 
        m82_1_1, N_83, bitalign_curr_state89, m23_1_2, 
        un1_bitalign_curr_state_14_1_Z, N_124_mux, m37_1_1, m37, 
        i12_mux_0, N_35, m7_1_1, N_8, tapcnt_final_2_sqmuxa, m86_1, 
        m85_1, N_76_0, m67_1, m66_1, N_51, N_119_mux, m55_0, 
        tapcnt_final_13_m0s2_0, un1_tapcnt_final_0_sqmuxa_Z, N_15, 
        m50_1_1, N_47, N_50, N_9, N_11, early_cur_set_0_sqmuxa_1_Z, 
        tapcnt_final_5_sqmuxa, rx_err_1_sqmuxa_Z, 
        calc_done_4_sqmuxa_0_Z, un1_bitalign_curr_state_0_sqmuxa_9_4_Z, 
        un1_bitalign_curr_state_0_sqmuxa_9_i, calc_done25_248, 
        calc_done25_249, calc_done25_168, calc_done25_169, 
        calc_done25_235, calc_done25_213, un34lto7_3, 
        tap_cnt_0_sqmuxa_0_Z, rx_BIT_ALGN_ERR_3_Z, reset_dly_fg4_4_Z, 
        early_late_diff_0_sqmuxa_1_0_Z, tap_cnt_0_sqmuxa_2_0, 
        un1_bitalign_curr_state_1_sqmuxa_2_i_0, N_63_0, 
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z, N_82, N_1498, N_1499, 
        un1_early_flags_pmux_1_Z, 
        un2_noearly_nolate_diff_start_validlt2, 
        bitalign_curr_state153_1_Z, bitalign_curr_state155_1, 
        bitalign_curr_state152_1_Z, un1_bitalign_curr_state_15_1_Z, 
        N_1416, un1_sig_re_train_Z, bitalign_curr_state149_1_Z, 
        bitalign_curr_state163_2, calc_done25_191, calc_done25_190, 
        calc_done25_189, calc_done25_188, calc_done25_187, 
        calc_done25_186, calc_done25_185, calc_done25_184, 
        calc_done25_183, calc_done25_182, calc_done25_181, 
        calc_done25_180, calc_done25_179, calc_done25_178, 
        calc_done25_177, calc_done25_176, calc_done25_175, 
        calc_done25_174, calc_done25_173, calc_done25_172, 
        calc_done25_171, calc_done25_170, calc_done25_167, 
        calc_done25_166, calc_done25_165, calc_done25_164, 
        calc_done25_163, calc_done25_162, calc_done25_161, 
        calc_done25_160, calc_done25_159, calc_done25_158, 
        calc_done25_157, calc_done25_156, calc_done25_155, 
        calc_done25_154, calc_done25_153, calc_done25_152, 
        calc_done25_151, calc_done25_150, calc_done25_149, 
        calc_done25_148, calc_done25_147, calc_done25_146, 
        calc_done25_145, calc_done25_144, calc_done25_143, 
        calc_done25_142, calc_done25_141, calc_done25_140, 
        calc_done25_139, calc_done25_138, calc_done25_137, 
        calc_done25_136, calc_done25_135, calc_done25_134, 
        calc_done25_133, calc_done25_132, calc_done25_131, 
        calc_done25_130, calc_done25_129, calc_done25_128, 
        bitalign_curr_state_2_sqmuxa_4_0_0, 
        un2_noearly_nolate_diff_nxt_validlto7_2_Z, 
        un2_noearly_nolate_diff_start_validlto7_2, 
        early_flags_dec_127_4_Z, un2_early_late_diff_validlto7_2_Z, 
        bit_align_dly_done_0_sqmuxa_1_0_Z, 
        rx_BIT_ALGN_MOVE_0_sqmuxa_0_Z, un34lto7_4, 
        tap_cnt_0_sqmuxa_1_0_Z, rx_BIT_ALGN_ERR_4_Z, reset_dly_fg4_6_Z, 
        un1_early_flags_1_sqmuxa_i, 
        un2_noearly_nolate_diff_nxt_validlt3, 
        bitalign_curr_state152_3_Z, un1_bitalign_curr_state151_Z, 
        bitalign_curr_state13, bitalign_curr_state61, N_114_mux, 
        bitalign_curr_state154_3_Z, N_31, 
        un1_bitalign_curr_state_16_1_Z, bitalign_curr_state12_0, 
        reset_dly_fg4_8_Z, bitalign_curr_state156_Z, 
        bitalign_curr_state153_Z, bitalign_curr_state161_Z, un34, 
        bitalign_curr_state155, bitalign_curr_state_0_sqmuxa_8_Z, 
        bitalign_curr_state163_Z, un2_early_late_diff_validlt7, 
        tapcnt_final_1_sqmuxa_2, N_61, un1_restart_trng_fg_0, N_108, 
        un1_bitalign_curr_state_1_sqmuxa_6_i_0, 
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z, 
        un1_bitalign_curr_state152_Z, bitalign_curr_state164_Z, 
        bitalign_curr_state154_Z, un1_calc_done25_7_i, 
        bitalign_curr_state61_0, bitalign_curr_state61_1_Z, 
        bitalign_curr_state61_4_Z, bitalign_curr_state61_5_Z, 
        bitalign_curr_state61_6_Z, bitalign_curr_state61_3_Z, 
        bitalign_curr_state61_2_Z, un1_bitalign_curr_state_15_0_Z, 
        calc_done25_231, calc_done25_230, calc_done25_229, 
        calc_done25_228, calc_done25_227, calc_done25_226, 
        calc_done25_225, calc_done25_224, 
        un1_bitalign_curr_state148_3_Z, un1_bitalign_curr_state148_2_Z, 
        rx_BIT_ALGN_LOAD_0_sqmuxa_Z, 
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_Z, N_52, CO1, 
        timeout_cnt_0_sqmuxa_Z, bit_align_done_0_sqmuxa_2_Z, N_98, 
        early_flags_1_sqmuxa_1_Z, emflag_cnt_0_sqmuxa_1_Z, 
        timeout_cnt_1_sqmuxa_Z, early_flags_0_sqmuxa_Z, 
        early_flags_1_sqmuxa_Z, rx_trng_done_1_sqmuxa_Z, 
        early_flags_0_sqmuxa_1_Z, bitalign_curr_state_1_sqmuxa_4_Z, 
        un1_rx_BIT_ALGN_LOAD_0_sqmuxa_i_0, N_14, 
        un1_bitalign_curr_state148_8_0_Z, 
        un1_bitalign_curr_state148_4_1_Z, 
        un1_bitalign_curr_state148_5_4_Z, 
        bitalign_curr_state_0_sqmuxa_9_Z, 
        bit_align_done_0_sqmuxa_3_1_Z, early_late_diff_0_sqmuxa_Z, 
        un1_noearly_nolate_diff_nxt_valid_Z, 
        un1_noearly_nolate_diff_start_valid, 
        un1_bitalign_curr_state148_8_1_Z, tapcnt_final_upd_3_sqmuxa_Z, 
        un1_early_flags_1_sqmuxa_1_Z, un1_bitalign_curr_state_13_1_Z, 
        bitalign_curr_state61_NE_4_Z, 
        un1_bitalign_curr_state_0_sqmuxa_9_1_Z, 
        un1_restart_trng_fg_10_0_Z, un1_bitalign_curr_state_15_2_Z, 
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_1_Z, 
        un1_bitalign_curr_state_14_1_0_Z, 
        un1_bitalign_curr_state148_5_Z, 
        un1_bitalign_curr_state_2_sqmuxa, emflag_cnt_1_sqmuxa_1_Z, 
        i22_mux, bitalign_curr_state_1_sqmuxa_7, 
        tapcnt_final_upd_2_sqmuxa, N_130_mux, emflag_cntlde_2, 
        un1_bitalign_curr_state148_8_2_Z, 
        un1_bitalign_curr_state148_9_2_Z, calc_done26, calc_done28, 
        un1_bitalign_curr_state_0_sqmuxa_9_2_Z;
    
    SLE \cnt[0]  (.D(CO0_0_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(CO0_0));
    SLE \early_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[4]));
    CFG3 #( .INIT(8'h40) )  rx_BIT_ALGN_MOVE_0_sqmuxa_0 (.A(
        bitalign_curr_state_Z[0]), .B(tap_cnt_0_sqmuxa_2_0), .C(
        bitalign_curr_state_Z[1]), .Y(rx_BIT_ALGN_MOVE_0_sqmuxa_0_Z));
    SLE \late_flags[59]  (.D(late_flags_7_fast_0[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[59]));
    SLE \early_flags[93]  (.D(early_flags_7_fast_0[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[93]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[46]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[46]), .C(
        un10_early_flags[46]), .Y(late_flags_7_fast_0[46]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_235  (.A(
        calc_done25_175), .B(calc_done25_174), .C(calc_done25_173), .D(
        calc_done25_172), .Y(calc_done25_235));
    SLE \late_flags[38]  (.D(late_flags_7_fast_0[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[38]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[27]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[27]), .C(
        un10_early_flags[27]), .Y(early_flags_7_fast_0[27]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_157  (.A(
        early_flags_Z[11]), .B(early_flags_Z[10]), .C(early_flags_Z[9])
        , .D(early_flags_Z[8]), .Y(calc_done25_157));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[125]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[125]), .C(
        un10_early_flags[125]), .Y(early_flags_7_fast_0[125]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_3 (.A(
        un10_early_flags_2_0[0]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[3]));
    CFG4 #( .INIT(16'h3332) )  \tapcnt_final_13_sn.m3  (.A(
        tapcnt_final_1_sqmuxa_2), .B(restart_trng_fg_i), .C(
        tapcnt_final_2_sqmuxa), .D(tapcnt_final_3_sqmuxa_Z), .Y(
        un1_bitalign_curr_state169_12_sn));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[87]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[87]), .C(
        un10_early_flags[87]), .Y(early_flags_7_fast_0[87]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[124]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[124]), .C(
        un10_early_flags[124]), .Y(early_flags_7_fast_0[124]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[61]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[61]), .C(
        un10_early_flags[61]), .Y(late_flags_7_fast_0[61]));
    SLE \early_flags[127]  (.D(early_flags_7_fast_0[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[127]));
    CFG4 #( .INIT(16'h0008) )  bitalign_curr_state12 (.A(
        reset_dly_fg_Z), .B(bitalign_curr_state12_0), .C(
        BIT_ALGN_ERR_c), .D(rx_trng_done_Z), .Y(
        bitalign_curr_state12_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_30 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[0]), .D(un10_early_flags_30_0_Z), .Y(
        un10_early_flags[30]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_10 (.A(
        late_flags_pmux_63_1_0_0_y21), .B(late_flags_pmux_63_1_0_0_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_63_1_0_co0_4), .S(
        late_flags_pmux_63_1_0_wmux_10_S_0), .Y(
        late_flags_pmux_63_1_0_wmux_10_Y_0), .FCO(
        late_flags_pmux_63_1_0_co1_4));
    SLE \late_flags[95]  (.D(late_flags_7_fast_0[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[95]));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_82 (.A(tap_cnt_Z[5]), 
        .B(N_1499), .C(un10_early_flags_2_Z[0]), .D(
        un10_early_flags_1_Z[64]), .Y(un10_early_flags[82]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[14]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[14]), .C(
        un10_early_flags[14]), .Y(late_flags_7_fast_0[14]));
    SLE \late_flags[24]  (.D(late_flags_7_fast_0[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[24]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_172  (.A(
        late_flags_Z[63]), .B(late_flags_Z[62]), .C(late_flags_Z[61]), 
        .D(late_flags_Z[60]), .Y(calc_done25_172));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_16 (.A(
        early_flags_pmux_126_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[45]), .D(early_flags_Z[109]), .FCI(
        early_flags_pmux_126_1_1_co0_7), .S(
        early_flags_pmux_126_1_1_wmux_16_S_0), .Y(
        early_flags_pmux_126_1_1_y5_0), .FCO(
        early_flags_pmux_126_1_1_co1_7));
    CFG2 #( .INIT(4'hB) )  rx_trng_done1_1_sqmuxa_i (.A(N_61), .B(
        bitalign_curr_state148_Z), .Y(N_52));
    CFG4 #( .INIT(16'hFFFE) )  emflag_cnt_0_sqmuxa_1_RNIESLM (.A(
        emflag_cnt_0_sqmuxa), .B(tap_cnt_0_sqmuxa_1_Z), .C(
        restart_trng_fg_i), .D(emflag_cnt_0_sqmuxa_1_Z), .Y(
        emflag_cntlde_2));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[82]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[82]), .C(
        un10_early_flags[82]), .Y(late_flags_7_fast_0[82]));
    SLE \late_flags[6]  (.D(late_flags_7_fast_0[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[67]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[67]), .C(
        un10_early_flags[67]), .Y(early_flags_7_fast_0[67]));
    CFG3 #( .INIT(8'h01) )  bitalign_curr_state41 (.A(wait_cnt_Z[2]), 
        .B(wait_cnt_Z[1]), .C(wait_cnt_Z[0]), .Y(
        bitalign_curr_state41_Z));
    SLE \noearly_nolate_diff_start[7]  (.D(
        noearly_nolate_diff_start_7[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_7));
    CFG4 #( .INIT(16'h0C5C) )  \bitalign_curr_state_34_4_0_.m62  (.A(
        N_35), .B(N_60_0), .C(bitalign_curr_state_Z[0]), .D(
        early_flags_dec[127]), .Y(N_63));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_2 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[0]), .D(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[2]));
    SLE rx_trng_done1 (.D(N_1415_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_trng_done1_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_trng_done1_Z));
    CFG3 #( .INIT(8'hFB) )  bit_align_dly_done_0_sqmuxa_1_i (.A(
        tap_cnt_0_sqmuxa_1_Z), .B(bit_align_done_0_sqmuxa_3_1_Z), .C(
        bitalign_curr_state_0_sqmuxa_9_Z), .Y(
        bit_align_dly_done_0_sqmuxa_1_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[92]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[92]), .C(
        un10_early_flags[92]), .Y(early_flags_7_fast_0[92]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_20 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[16]), .C(
        un10_early_flags_1_Z[20]), .Y(un10_early_flags[20]));
    SLE \late_flags[69]  (.D(late_flags_7_fast_0[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[69]));
    CFG4 #( .INIT(16'h5540) )  early_val_2_sqmuxa (.A(
        restart_trng_fg_i), .B(un1_early_last_set_1_sqmuxa_1_1_tz_Z), 
        .C(early_flags_pmux), .D(early_last_set_1_sqmuxa_1_3_Z), .Y(
        early_val_2_sqmuxa_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_0 (.A(
        late_flags_pmux_63_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[34]), .D(late_flags_Z[98]), .FCI(
        late_flags_pmux_63_1_0_0_co0), .S(
        late_flags_pmux_63_1_0_wmux_0_S_0), .Y(
        late_flags_pmux_63_1_0_0_y1), .FCO(
        late_flags_pmux_63_1_0_0_co1));
    SLE rx_BIT_ALGN_LOAD (.D(rx_BIT_ALGN_LOAD_9), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_BIT_ALGN_LOAD_0_sqmuxa_1_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD));
    SLE \late_flags[125]  (.D(late_flags_7_fast_0[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[125]));
    SLE \early_late_diff[1]  (.D(early_late_diff_8[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[1]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNIB02G2[4]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[4]), .D(GND), .FCI(
        timeout_cnt_cry[3]), .S(timeout_cnt_s[4]), .Y(
        timeout_cnt_RNIB02G2_Y_0[4]), .FCO(timeout_cnt_cry[4]));
    CFG4 #( .INIT(16'h0010) )  bitalign_curr_state153 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state153_1_Z), .D(bitalign_curr_state_Z[1]), .Y(
        bitalign_curr_state153_Z));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_6 (.A(
        un10_tapcnt_final_6), .B(un16_tapcnt_final_6), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_5_Z), .S(
        un10_tapcnt_final_cry_6_S_0), .Y(un10_tapcnt_final_cry_6_Y_0), 
        .FCO(un10_tapcnt_final_cry_6_Z));
    SLE \late_flags[74]  (.D(late_flags_7_fast_0[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[74]));
    CFG4 #( .INIT(16'hFFFE) )  emflag_cnt_1_sqmuxa_1_RNI2CFH1 (.A(
        bitalign_curr_state_1_sqmuxa_4_Z), .B(emflag_cnt_1_sqmuxa_1_Z), 
        .C(rx_err_1_sqmuxa_Z), .D(emflag_cntlde_2), .Y(emflag_cnte));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_94 (.A(tap_cnt_Z[5]), 
        .B(un10_early_flags_1_Z[6]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[64]), .Y(un10_early_flags[94]));
    SLE \early_flags[34]  (.D(early_flags_7_fast_0[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[34]));
    CFG4 #( .INIT(16'hF800) )  un1_noearly_nolate_diff_nxt_valid (.A(
        un16_tapcnt_final_3), .B(un2_noearly_nolate_diff_nxt_validlt3), 
        .C(un2_noearly_nolate_diff_nxt_validlto7_2_Z), .D(
        un1_early_late_diff_1_cry_7_Z), .Y(
        un1_noearly_nolate_diff_nxt_valid_Z));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNIEOFU2[5]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[5]), .D(GND), .FCI(
        timeout_cnt_cry[4]), .S(timeout_cnt_s[5]), .Y(
        timeout_cnt_RNIEOFU2_Y_0[5]), .FCO(timeout_cnt_cry[5]));
    SLE \early_flags[40]  (.D(early_flags_7_fast_0[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[40]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[108]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[108]), .C(
        un10_early_flags[108]), .Y(late_flags_7_fast_0[108]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_9_1 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[9]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[31]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[31]), .C(
        un10_early_flags[31]), .Y(early_flags_7_fast_0[31]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[12]), 
        .D(late_flags_Z[76]), .FCI(late_flags_pmux_63_1_1_co1_6), .S(
        late_flags_pmux_63_1_1_wmux_15_S_0), .Y(
        late_flags_pmux_63_1_1_y0_6), .FCO(
        late_flags_pmux_63_1_1_co0_7));
    SLE \early_flags[5]  (.D(early_flags_7_fast_0[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[5]));
    SLE \late_flags[34]  (.D(late_flags_7_fast_0[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[34]));
    SLE \late_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[2])
        );
    SLE \timeout_cnt[7]  (.D(timeout_cnt_s[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[7]));
    SLE \restart_reg[2]  (.D(restart_reg_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_reg_Z[2]));
    SLE \early_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[5]));
    SLE \no_early_no_late_val_st2[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[2]));
    SLE \tapcnt_final_upd[1]  (.D(tapcnt_final_upd_8_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[1]));
    SLE \noearly_nolate_diff_nxt[7]  (.D(noearly_nolate_diff_nxt_8[7]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_7));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[26]), 
        .D(early_flags_Z[90]), .FCI(early_flags_pmux_63_1_0_co1_1), .S(
        early_flags_pmux_63_1_0_wmux_5_S_0), .Y(
        early_flags_pmux_63_1_0_y0_2), .FCO(
        early_flags_pmux_63_1_0_co0_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[29]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[29]), .C(
        un10_early_flags[29]), .Y(early_flags_7_fast_0[29]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[8]), .D(
        late_flags_Z[72]), .FCI(late_flags_pmux_63_1_1_co1_0), .S(
        late_flags_pmux_63_1_1_wmux_3_S_0), .Y(
        late_flags_pmux_63_1_1_y0_1), .FCO(
        late_flags_pmux_63_1_1_co0_1));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_111_1_0 (.A(
        un10_early_flags_1_Z[3]), .B(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags_1_0[15]));
    CFG4 #( .INIT(16'hAAAB) )  rx_BIT_ALGN_DIR_0_sqmuxa_2_i (.A(
        restart_trng_fg_i), .B(un1_bitalign_curr_state_15_2_Z), .C(
        early_flags_0_sqmuxa_1_Z), .D(tapcnt_final_upd_3_sqmuxa_Z), .Y(
        rx_BIT_ALGN_DIR_0_sqmuxa_2_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[89]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[89]), .C(
        un10_early_flags[89]), .Y(early_flags_7_fast_0[89]));
    SLE \early_flags[64]  (.D(early_flags_7_fast_0[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[64]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[22]), 
        .D(early_flags_Z[86]), .FCI(early_flags_pmux_63_1_0_co1_5), .S(
        early_flags_pmux_63_1_0_wmux_13_S_0), .Y(
        early_flags_pmux_63_1_0_y0_5), .FCO(
        early_flags_pmux_63_1_0_co0_6));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_249  (.A(
        calc_done25_231), .B(calc_done25_230), .C(calc_done25_229), .D(
        calc_done25_228), .Y(calc_done25_249));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_5 (.A(late_val_Z[5])
        , .B(early_val_Z[5]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_4_Z), .S(tapcnt_final27_cry_5_S_0), .Y(
        tapcnt_final27_cry_5_Y_0), .FCO(tapcnt_final27_cry_5_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_13_1 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[5]));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[2]  (.A(
        tapcnt_final_13_Z[3]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[2]), .Y(tapcnt_final_13_1_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[63]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[63]), .C(
        un10_early_flags[63]), .Y(late_flags_7_fast_0[63]));
    CFG4 #( .INIT(16'hFFA8) )  
        \bitalign_curr_state_34_4_0_.un2_noearly_nolate_diff_start_validlto7  
        (.A(un10_tapcnt_final_3), .B(un10_tapcnt_final_2), .C(
        un2_noearly_nolate_diff_start_validlt2), .D(
        un2_noearly_nolate_diff_start_validlto7_2), .Y(
        un2_noearly_nolate_diff_start_valid));
    CFG2 #( .INIT(4'hE) )  un1_restart_trng_fg_10_1 (.A(
        bitalign_curr_state_1_sqmuxa_4_Z), .B(restart_trng_fg_i), .Y(
        un1_restart_trng_fg_10_sn_1));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[3]  (.A(
        tapcnt_final_13_Z[4]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[3]), .Y(tapcnt_final_13_1_Z[3]));
    SLE \early_flags[36]  (.D(early_flags_7_fast_0[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[36]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[114]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[114]), .C(
        un10_early_flags[114]), .Y(late_flags_7_fast_0[114]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_147  (.A(
        early_flags_Z[59]), .B(early_flags_Z[58]), .C(
        early_flags_Z[57]), .D(early_flags_Z[56]), .Y(calc_done25_147));
    SLE \late_flags[110]  (.D(late_flags_7_fast_0[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[110]));
    SLE \early_flags[37]  (.D(early_flags_7_fast_0[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[37]));
    SLE \early_flags[105]  (.D(early_flags_7_fast_0[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[105]));
    SLE \early_flags[118]  (.D(early_flags_7_fast_0[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[118]));
    CFG3 #( .INIT(8'hE4) )  \early_flags_RNO[49]  (.A(N_208), .B(
        EYE_MONITOR_EARLY_net_0_0), .C(early_flags_Z[49]), .Y(
        early_flags_RNO_0[49]));
    CFG2 #( .INIT(4'hE) )  un1_restart_trng_fg_5 (.A(
        un1_tap_cnt_0_sqmuxa_6_0), .B(restart_trng_fg_i), .Y(
        un1_restart_trng_fg_5_0));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_12 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[12]));
    SLE \early_flags[120]  (.D(early_flags_7_fast_0[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[120]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[69]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[69]), .C(
        un10_early_flags[69]), .Y(early_flags_7_fast_0[69]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_12 (.A(
        late_flags_pmux_63_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[38]), .D(late_flags_Z[102]), .FCI(
        late_flags_pmux_63_1_0_co0_5), .S(
        late_flags_pmux_63_1_0_wmux_12_S_0), .Y(
        late_flags_pmux_63_1_0_y1_0), .FCO(
        late_flags_pmux_63_1_0_co1_5));
    SLE \early_flags[31]  (.D(early_flags_7_fast_0[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[31]));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_46_3 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_3_Z[46]));
    SLE \early_flags[15]  (.D(early_flags_7_fast_0[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[15]));
    CFG4 #( .INIT(16'h7FFF) )  
        \bitalign_curr_state_34_4_0_.calc_done25_253_1_0  (.A(
        calc_done25_239), .B(calc_done25_238), .C(calc_done25_233), .D(
        calc_done25_232), .Y(calc_done25_253_1_0));
    SLE \early_flags[42]  (.D(early_flags_7_fast_0[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[42]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_85 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[5]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[4]), .Y(
        un10_early_flags[85]));
    CFG4 #( .INIT(16'h7340) )  \bitalign_curr_state_34_4_0_.m40_1_1  (
        .A(bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[4]), .C(
        N_124_mux), .D(N_15), .Y(m40_1_1));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_161  (.A(
        late_flags_Z[11]), .B(late_flags_Z[10]), .C(late_flags_Z[9]), 
        .D(late_flags_Z[8]), .Y(calc_done25_161));
    SLE \noearly_nolate_diff_nxt[1]  (.D(noearly_nolate_diff_nxt_8[1]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_1));
    SLE \no_early_no_late_val_end2[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[5]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[5]), .C(
        un10_early_flags[5]), .Y(late_flags_7_fast_0[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[2]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[2]), .C(
        un10_early_flags[2]), .Y(late_flags_7_fast_0[2]));
    SLE \early_flags[66]  (.D(early_flags_7_fast_0[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[66]));
    CFG4 #( .INIT(16'hFFFE) )  restart_trng_fg (.A(
        restart_edge_reg_Z[3]), .B(restart_edge_reg_Z[2]), .C(
        restart_edge_reg_Z[1]), .D(restart_edge_reg_Z[0]), .Y(
        restart_trng_fg_i));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_14 (.A(
        early_flags_pmux_126_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[53]), .D(early_flags_Z[117]), .FCI(
        early_flags_pmux_126_1_1_co0_6), .S(
        early_flags_pmux_126_1_1_wmux_14_S_0), .Y(
        early_flags_pmux_126_1_1_y3_0), .FCO(
        early_flags_pmux_126_1_1_co1_6));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.m43_0_a2  (.A(
        bitalign_curr_state12_Z), .B(un1_rx_BIT_ALGN_START), .Y(
        bitalign_curr_state13));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_189  (.A(
        late_flags_Z[99]), .B(late_flags_Z[98]), .C(late_flags_Z[97]), 
        .D(late_flags_Z[96]), .Y(calc_done25_189));
    SLE \early_flags[67]  (.D(early_flags_7_fast_0[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[67]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_2 (.A(
        early_flags_pmux_63_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[48]), .D(early_flags_Z[112]), .FCI(
        early_flags_pmux_63_1_1_co0_0), .S(
        early_flags_pmux_63_1_1_wmux_2_S_0), .Y(
        early_flags_pmux_63_1_1_y3), .FCO(
        early_flags_pmux_63_1_1_co1_0));
    SLE \early_flags[74]  (.D(early_flags_7_fast_0[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[74]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[92]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[92]), .C(
        un10_early_flags[92]), .Y(late_flags_7_fast_0[92]));
    SLE \early_flags[119]  (.D(early_flags_7_fast_0[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[119]));
    SLE \early_flags[61]  (.D(early_flags_7_fast_0[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[61]));
    SLE \timeout_cnt[4]  (.D(timeout_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[84]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[84]), .C(
        un10_early_flags[84]), .Y(late_flags_7_fast_0[84]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[122]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[122]), .C(
        un10_early_flags[122]), .Y(early_flags_7_fast_0[122]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_32_1_0_a2 (.A(tap_cnt_Z[5])
        , .B(tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[32]));
    SLE \wait_cnt[2]  (.D(wait_cnt_4_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(wait_cnt_Z[2]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_4_0 (
        .A(emflag_cnt_Z[4]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[4]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_3), .S(
        noearly_nolate_diff_start_7[4]), .Y(
        noearly_nolate_diff_start_7_cry_4_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_4));
    CFG4 #( .INIT(16'h53FF) )  \bitalign_curr_state_34_4_0_.m64_1_1  (
        .A(bitalign_curr_state41_Z), .B(N_60_0), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        m64_1_1));
    CFG1 #( .INIT(2'h1) )  un1_restart_trng_fg_5_RNIIB4C (.A(
        un1_restart_trng_fg_5_0), .Y(N_19_i));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_126 (.A(tap_cnt_Z[0]), 
        .B(un10_early_flags_1_Z[6]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[126]));
    SLE \late_flags[82]  (.D(late_flags_7_fast_0[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[82]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_59 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_2_Z[35]), .Y(
        un10_early_flags[59]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_35_2 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[35]));
    SLE \noearly_nolate_diff_nxt[0]  (.D(noearly_nolate_diff_nxt_8[0]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_0));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[113]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[113]), .C(
        un10_early_flags[113]), .Y(late_flags_7_fast_0[113]));
    SLE \late_flags[102]  (.D(late_flags_7_fast_0[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[102]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_87_3 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_3_Z[87]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[106]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[106]), .C(
        un10_early_flags[106]), .Y(late_flags_7_fast_0[106]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[97]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[97]), .C(
        un10_early_flags[97]), .Y(early_flags_7_fast_0[97]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[14]), 
        .D(early_flags_Z[78]), .FCI(early_flags_pmux_63_1_0_co1_6), .S(
        early_flags_pmux_63_1_0_wmux_15_S_0), .Y(
        early_flags_pmux_63_1_0_y0_6), .FCO(
        early_flags_pmux_63_1_0_co0_7));
    CFG4 #( .INIT(16'h0020) )  bit_align_done_2_sqmuxa (.A(
        bit_align_dly_done_0_sqmuxa_1_0_Z), .B(restart_trng_fg_i), .C(
        bitalign_curr_state161_2_Z), .D(sig_re_train_Z), .Y(
        bit_align_done_2_sqmuxa_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_131  (.A(
        early_flags_Z[123]), .B(early_flags_Z[122]), .C(
        early_flags_Z[121]), .D(early_flags_Z[120]), .Y(
        calc_done25_131));
    CFG4 #( .INIT(16'h00E0) )  sig_re_train (.A(
        EYE_MONITOR_LATE_net_0_0), .B(EYE_MONITOR_EARLY_net_0_0), .C(
        un1_sig_re_train_Z), .D(BIT_ALGN_ERR_c), .Y(sig_re_train_Z));
    SLE \late_flags[12]  (.D(late_flags_7_fast_0[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[12]));
    SLE \early_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[3]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_69 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[64]), .C(
        un10_early_flags_2_Z[69]), .Y(un10_early_flags[69]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_14 (.A(
        early_flags_pmux_126_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[55]), .D(early_flags_Z[119]), .FCI(
        early_flags_pmux_126_1_0_co0_6), .S(
        early_flags_pmux_126_1_0_wmux_14_S_0), .Y(
        early_flags_pmux_126_1_0_y3_0), .FCO(
        early_flags_pmux_126_1_0_co1_6));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_117 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_1_Z[48]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_2_Z[69]), .Y(
        un10_early_flags[117]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[56]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[56]), .C(
        un10_early_flags[56]), .Y(early_flags_7_fast_0[56]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[72]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[72]), .C(
        un10_early_flags[72]), .Y(early_flags_7_fast_0[72]));
    SLE \early_flags[76]  (.D(early_flags_7_fast_0[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[76]));
    CFG4 #( .INIT(16'h0FEE) )  \bitalign_curr_state_34_4_0_.m82_1_0  (
        .A(BIT_ALGN_ERR_c), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .C(N_63), 
        .D(bitalign_curr_state_Z[1]), .Y(m82_1_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[18]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[18]), .C(
        un10_early_flags[18]), .Y(early_flags_7_fast_0[18]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_97 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_2_Z[69]), .D(
        un10_early_flags_2_0[96]), .Y(un10_early_flags[97]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_34 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_2_0[32]), .Y(un10_early_flags[34]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[10]), 
        .D(early_flags_Z[74]), .FCI(early_flags_pmux_63_1_0_co1_0), .S(
        early_flags_pmux_63_1_0_wmux_3_S_0), .Y(
        early_flags_pmux_63_1_0_y0_1), .FCO(
        early_flags_pmux_63_1_0_co0_1));
    SLE \early_flags[77]  (.D(early_flags_7_fast_0[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[77]));
    SLE \no_early_no_late_val_end1[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[4]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_88 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_1_Z[64]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[88]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_14 (.A(
        early_flags_pmux_63_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[54]), .D(early_flags_Z[118]), .FCI(
        early_flags_pmux_63_1_0_co0_6), .S(
        early_flags_pmux_63_1_0_wmux_14_S_0), .Y(
        early_flags_pmux_63_1_0_y3_0), .FCO(
        early_flags_pmux_63_1_0_co1_6));
    SLE \early_flags[111]  (.D(early_flags_7_fast_0[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[111]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_37_2_0_a2 (.A(tap_cnt_Z[5])
        , .B(tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[37]));
    SLE \late_flags[42]  (.D(late_flags_7_fast_0[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[42]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[15]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[15]), .C(
        un10_early_flags[15]), .Y(early_flags_7_fast_0[15]));
    SLE \early_flags[71]  (.D(early_flags_7_fast_0[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[71]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[69]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[69]), .C(
        un10_early_flags[69]), .Y(late_flags_7_fast_0[69]));
    CFG4 #( .INIT(16'hFFFE) )  rx_BIT_ALGN_LOAD_0_sqmuxa_1_i (.A(
        restart_trng_fg_i), .B(rx_BIT_ALGN_LOAD_0_sqmuxa_Z), .C(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .D(
        un1_tap_cnt_0_sqmuxa_6_0), .Y(rx_BIT_ALGN_LOAD_0_sqmuxa_1_i_Z));
    SLE \bitalign_curr_state[4]  (.D(bitalign_curr_state_34[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[4]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_19 (.A(
        early_flags_pmux_126_1_0_y7_0), .B(
        early_flags_pmux_126_1_0_y5_0), .C(emflag_cnt_Z[4]), .D(
        emflag_cnt_Z[3]), .FCI(early_flags_pmux_126_1_0_co1_8), .S(
        early_flags_pmux_126_1_0_wmux_19_S_0), .Y(
        early_flags_pmux_126_1_0_y0_8), .FCO(
        early_flags_pmux_126_1_0_co0_9));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[113]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[113]), .C(
        un10_early_flags[113]), .Y(early_flags_7_fast_0[113]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_19 (.A(
        late_flags_pmux_126_1_0_y7_0), .B(late_flags_pmux_126_1_0_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co1_8), .S(
        late_flags_pmux_126_1_0_wmux_19_S_0), .Y(
        late_flags_pmux_126_1_0_y0_8), .FCO(
        late_flags_pmux_126_1_0_co0_9));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_119 (.A(
        un10_early_flags_1_Z[20]), .B(tap_cnt_Z[3]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[96]), .Y(
        un10_early_flags[119]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_7 (.A(
        late_flags_pmux_126_1_0_0_y7), .B(late_flags_pmux_126_1_0_0_y5)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co1_2), .S(
        late_flags_pmux_126_1_0_wmux_7_S_0), .Y(
        late_flags_pmux_126_1_0_y0_3), .FCO(
        late_flags_pmux_126_1_0_co0_3));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_163  (.A(
        late_flags_Z[3]), .B(late_flags_Z[2]), .C(late_flags_Z[1]), .D(
        late_flags_Z[0]), .Y(calc_done25_163));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_24 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_2_0[24]), .C(
        un10_early_flags_1_Z[0]), .Y(un10_early_flags[24]));
    SLE \early_flags[113]  (.D(early_flags_7_fast_0[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[113]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_2_0 (
        .A(emflag_cnt_Z[2]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[2]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_1), .S(
        noearly_nolate_diff_start_7[2]), .Y(
        noearly_nolate_diff_start_7_cry_2_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[46]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[46]), .C(
        un10_early_flags[46]), .Y(early_flags_7_fast_0[46]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_15 (.A(
        un10_early_flags_2_0[0]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[15]));
    CFG4 #( .INIT(16'h2232) )  \bitalign_curr_state_34_4_0_.m91_1  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        un1_retrain_adj_tap_i), .D(N_69), .Y(m91_1_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[121]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[121]), .C(
        un10_early_flags[121]), .Y(early_flags_7_fast_0[121]));
    SLE \timeout_cnt[3]  (.D(timeout_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[3]));
    CFG4 #( .INIT(16'h0008) )  
        \bitalign_curr_state_34_4_0_.calc_done27  (.A(
        un2_noearly_nolate_diff_start_valid), .B(
        un1_early_late_diff_cry_7_Z), .C(calc_done25), .D(
        un1_tapcnt_final), .Y(calc_done27));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_233  (.A(
        calc_done25_167), .B(calc_done25_166), .C(calc_done25_165), .D(
        calc_done25_164), .Y(calc_done25_233));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_18 (.A(
        early_flags_pmux_63_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[62]), .D(early_flags_Z[126]), .FCI(
        early_flags_pmux_63_1_0_co0_8), .S(
        early_flags_pmux_63_1_0_wmux_18_S_0), .Y(
        early_flags_pmux_63_1_0_y7_0), .FCO(
        early_flags_pmux_63_1_0_co1_8));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[0]  (.A(
        un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_Y_0[0]), .B(N_63_0), .Y(
        N_32_i));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_107 (.A(
        un10_early_flags_1_Z[40]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_2_Z[67]), .Y(
        un10_early_flags[107]));
    SLE \timeout_cnt[1]  (.D(timeout_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[1]));
    SLE \early_flags[38]  (.D(early_flags_7_fast_0[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[38]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_96 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_1_Z[96]), .C(
        un10_early_flags_2_0[96]), .Y(un10_early_flags[96]));
    SLE \late_flags[113]  (.D(late_flags_7_fast_0[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[113]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[1]), .D(
        late_flags_Z[65]), .FCI(VCC), .S(
        late_flags_pmux_126_1_1_wmux_S_0), .Y(
        late_flags_pmux_126_1_1_y0), .FCO(late_flags_pmux_126_1_1_co0));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[31]), 
        .D(early_flags_Z[95]), .FCI(early_flags_pmux_126_1_0_co1_7), 
        .S(early_flags_pmux_126_1_0_wmux_17_S_0), .Y(
        early_flags_pmux_126_1_0_y0_7), .FCO(
        early_flags_pmux_126_1_0_co0_8));
    SLE \retrain_reg[0]  (.D(sig_re_train_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(retrain_reg_Z[0]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[3]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[3]), .D(GND), .FCI(
        emflag_cnt_cry_Z[2]), .S(emflag_cnt_s[3]), .Y(
        emflag_cnt_cry_Y_1[3]), .FCO(emflag_cnt_cry_Z[3]));
    CFG4 #( .INIT(16'h0400) )  bitalign_curr_state154_3 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[2]), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state154_3_Z));
    SLE \restart_edge_reg[2]  (.D(restart_edge_reg_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[2]));
    CFG4 #( .INIT(16'h8000) )  reset_dly_fg4_6 (.A(rst_cnt_Z[5]), .B(
        rst_cnt_Z[4]), .C(rst_cnt_Z[3]), .D(rst_cnt_Z[2]), .Y(
        reset_dly_fg4_6_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[21]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[21]), .C(
        un10_early_flags[21]), .Y(early_flags_7_fast_0[21]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_40_1 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_1_Z[40]));
    SLE \early_flags[29]  (.D(early_flags_7_fast_0[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[29]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[81]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[81]), .C(
        un10_early_flags[81]), .Y(early_flags_7_fast_0[81]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_162  (.A(
        late_flags_Z[7]), .B(late_flags_Z[6]), .C(late_flags_Z[5]), .D(
        late_flags_Z[4]), .Y(calc_done25_162));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIJGIR[1]  (.A(
        late_val_Z[1]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[1]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIJGIR_0[1]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[99]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[99]), .C(
        un10_early_flags[99]), .Y(early_flags_7_fast_0[99]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[66]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[66]), .C(
        un10_early_flags[66]), .Y(late_flags_7_fast_0[66]));
    CFG2 #( .INIT(4'h2) )  Restart_trng_edge_det (.A(restart_reg_Z[1]), 
        .B(restart_reg_Z[2]), .Y(Restart_trng_edge_det_Z));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_81 (.A(N_1498), .B(
        tap_cnt_Z[5]), .C(un10_early_flags_2_Z[69]), .D(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[81]));
    CFG4 #( .INIT(16'h00AC) )  \bitalign_curr_state_34_4_0_.m41  (.A(
        N_40), .B(m40_1_1), .C(bitalign_curr_state_Z[3]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[0]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_1_wmux_20 (.A(
        late_flags_pmux_63_1_1_y0_8), .B(late_flags_pmux_63_1_1_y3_0), 
        .C(late_flags_pmux_63_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co0_9), .S(
        late_flags_pmux_63_1_1_wmux_20_S_0), .Y(
        late_flags_pmux_63_1_1_y21), .FCO(late_flags_pmux_63_1_1_co1_9)
        );
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_0 (.A(
        un10_tapcnt_final_0), .B(early_late_diff_Z[0]), .C(GND), .D(
        GND), .FCI(GND), .S(un1_early_late_diff_cry_0_S_0), .Y(
        un1_early_late_diff_cry_0_Y_0), .FCO(
        un1_early_late_diff_cry_0_Z));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_109 (.A(
        un10_early_flags_2_Z[69]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[5]), .D(un10_early_flags_1_Z[40]), .Y(
        un10_early_flags[109]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_2 (.A(late_val_Z[2])
        , .B(early_val_Z[2]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_1_Z), .S(tapcnt_final27_cry_2_S_0), .Y(
        tapcnt_final27_cry_2_Y_0), .FCO(tapcnt_final27_cry_2_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_133  (.A(
        early_flags_Z[99]), .B(early_flags_Z[98]), .C(
        early_flags_Z[97]), .D(early_flags_Z[96]), .Y(calc_done25_133));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_12_1 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[12]));
    CFG2 #( .INIT(4'h2) )  late_last_set15 (.A(early_last_set_Z), .B(
        late_last_set_Z), .Y(late_last_set15_Z));
    SLE \late_flags[111]  (.D(late_flags_7_fast_0[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[111]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNIT5J81[0]  (.A(early_val_Z[0])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[0]), .Y(
        early_val_RNIT5J81_Z[0]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNO[7]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[7]), .D(GND), .FCI(
        timeout_cnt_cry[6]), .S(timeout_cnt_s[7]), .Y(
        timeout_cnt_RNO_Y_0[7]), .FCO(timeout_cnt_RNO_FCO_0[7]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_12 (.A(
        early_flags_pmux_126_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[37]), .D(early_flags_Z[101]), .FCI(
        early_flags_pmux_126_1_1_co0_5), .S(
        early_flags_pmux_126_1_1_wmux_12_S_0), .Y(
        early_flags_pmux_126_1_1_y1_0), .FCO(
        early_flags_pmux_126_1_1_co1_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[126]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[126]), .C(
        un10_early_flags[126]), .Y(late_flags_7_fast_0[126]));
    CFG2 #( .INIT(4'h8) )  calc_done_4_sqmuxa_0 (.A(
        bitalign_curr_state162_Z), .B(un1_early_late_diff_valid_Z), .Y(
        calc_done_4_sqmuxa_0_Z));
    SLE \late_flags[92]  (.D(late_flags_7_fast_0[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[92]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[61]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[61]), .C(
        un10_early_flags[61]), .Y(early_flags_7_fast_0[61]));
    SLE \early_flags[68]  (.D(early_flags_7_fast_0[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[68]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_11_1 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_1_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[94]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[94]), .C(
        un10_early_flags[94]), .Y(late_flags_7_fast_0[94]));
    SLE \bitalign_curr_state[0]  (.D(bitalign_curr_state_34[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[0]));
    CFG2 #( .INIT(4'h8) )  bitalign_curr_state152_1 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[1]), .Y(
        bitalign_curr_state152_1_Z));
    CFG2 #( .INIT(4'h2) )  rx_BIT_ALGN_START (.A(bit_align_start_Z), 
        .B(BIT_ALGN_ERR_c), .Y(BIT_ALGN_START_0_c));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[51]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[51]), .C(
        un10_early_flags[51]), .Y(late_flags_7_fast_0[51]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIBEUF3[0]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIHEIR_0[0]), .B(
        early_val_RNIT5J81_Z[0]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[0]), .FCI(GND), .S(early_val_RNIBEUF3_S[0]), .Y(
        early_val_RNIBEUF3_Y[0]), .FCO(tapcnt_final_13_m1_cry_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[0]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[0]), .C(
        un10_early_flags[0]), .Y(early_flags_7_fast_0[0]));
    CFG4 #( .INIT(16'h0F1B) )  \bitalign_curr_state_34_4_0_.m23  (.A(
        early_flags_dec[127]), .B(m23_1_2), .C(
        bitalign_curr_state_Z[1]), .D(un1_bitalign_curr_state_14_1_Z), 
        .Y(N_124_mux));
    CFG3 #( .INIT(8'h40) )  un10_early_flags_18 (.A(N_1499), .B(
        un10_early_flags_2_Z[10]), .C(un10_early_flags_2_0[16]), .Y(
        un10_early_flags[18]));
    CFG4 #( .INIT(16'hEFEE) )  un1_bitalign_curr_state_0_sqmuxa_9_1 (
        .A(early_flags_0_sqmuxa_Z), .B(
        bitalign_curr_state_0_sqmuxa_8_Z), .C(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .D(bitalign_curr_state154_Z), 
        .Y(un1_bitalign_curr_state_0_sqmuxa_9_1_Z));
    CFG4 #( .INIT(16'hFFFE) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i (
        .A(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .B(
        un1_bitalign_curr_state_1_sqmuxa_6_i_0), .C(restart_trng_fg_i), 
        .D(un1_rx_BIT_ALGN_LOAD_0_sqmuxa_i_0), .Y(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i_Z));
    SLE \late_flags[56]  (.D(late_flags_7_fast_0[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[56]));
    SLE \early_flags[102]  (.D(early_flags_7_fast_0[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[102]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_132  (.A(
        early_flags_Z[103]), .B(early_flags_Z[102]), .C(
        early_flags_Z[101]), .D(early_flags_Z[100]), .Y(
        calc_done25_132));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_2 (.A(
        late_flags_pmux_63_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[48]), .D(late_flags_Z[112]), .FCI(
        late_flags_pmux_63_1_1_co0_0), .S(
        late_flags_pmux_63_1_1_wmux_2_S_0), .Y(
        late_flags_pmux_63_1_1_y3), .FCO(late_flags_pmux_63_1_1_co1_0));
    SLE \late_flags[20]  (.D(late_flags_7_fast_0[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[20]));
    CFG3 #( .INIT(8'h20) )  early_last_set_1_sqmuxa_1_3 (.A(N_20), .B(
        late_last_set15_Z), .C(bitalign_curr_state161_Z), .Y(
        early_last_set_1_sqmuxa_1_3_Z));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_1_wmux_20 (.A(
        early_flags_pmux_126_1_1_y0_8), .B(
        early_flags_pmux_126_1_1_y3_0), .C(
        early_flags_pmux_126_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_1_co0_9), .S(
        early_flags_pmux_126_1_1_wmux_20_S_0), .Y(
        early_flags_pmux_126_1_1_y21), .FCO(
        early_flags_pmux_126_1_1_co1_9));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_8 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[3]), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[8]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[127]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[127]), .C(
        un10_early_flags[127]), .Y(early_flags_7_fast_0[127]));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_80 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[0]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[0]), .Y(
        un10_early_flags[80]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_1_0 (.A(
        emflag_cnt_Z[1]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[1]), .D(GND), .FCI(early_late_diff_8_cry_0), .S(
        early_late_diff_8[1]), .Y(early_late_diff_8_cry_1_0_Y_0), .FCO(
        early_late_diff_8_cry_1));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_2 (.A(
        un16_tapcnt_final_2), .B(un10_tapcnt_final_2), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_1_Z), .S(
        un16_tapcnt_final_cry_2_S_0), .Y(un16_tapcnt_final_cry_2_Y_0), 
        .FCO(un16_tapcnt_final_cry_2_Z));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_245  (.A(
        calc_done25_168), .B(calc_done25_169), .C(calc_done25_235), .D(
        calc_done25_213), .Y(calc_done25_245));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_9 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_126_1_0_co1_3), .S(
        early_flags_pmux_126_1_0_wmux_9_S_0), .Y(
        early_flags_pmux_126_1_0_wmux_9_Y_0), .FCO(
        early_flags_pmux_126_1_0_co0_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[77]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[77]), .C(
        un10_early_flags[77]), .Y(early_flags_7_fast_0[77]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_2 (.A(
        late_flags_pmux_126_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[49]), .D(late_flags_Z[113]), .FCI(
        late_flags_pmux_126_1_1_co0_0), .S(
        late_flags_pmux_126_1_1_wmux_2_S_0), .Y(
        late_flags_pmux_126_1_1_y3), .FCO(
        late_flags_pmux_126_1_1_co1_0));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[109]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[109]), .C(
        un10_early_flags[109]), .Y(late_flags_7_fast_0[109]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[13]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[13]), .C(
        un10_early_flags[13]), .Y(early_flags_7_fast_0[13]));
    CFG4 #( .INIT(16'h08FF) )  un1_early_flags_pmux_1_RNI26QC (.A(
        late_last_set15_Z), .B(bitalign_curr_state161_Z), .C(
        un1_early_flags_pmux_1_Z), .D(early_late_diff_0_sqmuxa_1_0_Z), 
        .Y(no_early_no_late_val_end2_0_sqmuxa_i));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_37 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[32]), .C(
        un10_early_flags_2_Z[37]), .Y(un10_early_flags[37]));
    SLE \tap_cnt[6]  (.D(N_1496_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tap_cnt_Z[6]));
    CFG2 #( .INIT(4'hE) )  rx_BIT_ALGN_DONE (.A(bit_align_done_Z), .B(
        BIT_ALGN_ERR_c), .Y(BIT_ALGN_DONE_0_c));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_10 (.A(
        late_flags_pmux_126_1_0_0_y21), .B(
        late_flags_pmux_126_1_0_0_y9), .C(emflag_cnt_Z[2]), .D(VCC), 
        .FCI(late_flags_pmux_126_1_0_co0_4), .S(
        late_flags_pmux_126_1_0_wmux_10_S_0), .Y(
        late_flags_pmux_126_1_0_wmux_10_Y_0), .FCO(
        late_flags_pmux_126_1_0_co1_4));
    SLE \early_flags[78]  (.D(early_flags_7_fast_0[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[78]));
    CFG4 #( .INIT(16'h0200) )  tapcnt_final_upd_2_sqmuxa_0_a2 (.A(
        mv_up_fg_Z), .B(mv_dn_fg_Z), .C(bitalign_curr_state12_Z), .D(
        N_98), .Y(tapcnt_final_upd_2_sqmuxa));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_0 (.A(
        early_flags_pmux_63_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[34]), .D(early_flags_Z[98]), .FCI(
        early_flags_pmux_63_1_0_0_co0), .S(
        early_flags_pmux_63_1_0_wmux_0_S_0), .Y(
        early_flags_pmux_63_1_0_0_y1), .FCO(
        early_flags_pmux_63_1_0_0_co1));
    CFG4 #( .INIT(16'h3AFA) )  \bitalign_curr_state_34_4_0_.m67_1  (.A(
        N_51), .B(N_119_mux), .C(bitalign_curr_state_Z[4]), .D(m55_0), 
        .Y(m67_1));
    SLE \late_flags[70]  (.D(late_flags_7_fast_0[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[70]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_48_2_0 (.A(
        un10_early_flags_2_Z[0]), .B(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[48]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_3_0 (.A(
        emflag_cnt_Z[3]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[3]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_2), .S(
        noearly_nolate_diff_nxt_8[3]), .Y(
        noearly_nolate_diff_nxt_8_cry_3_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_3));
    SLE \noearly_nolate_diff_start[0]  (.D(
        noearly_nolate_diff_start_7[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_0));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_42 (.A(
        un10_early_flags_1_Z[10]), .B(un10_early_flags_1_Z[32]), .C(
        un10_early_flags_2_0[40]), .Y(un10_early_flags[42]));
    CFG3 #( .INIT(8'hFD) )  rx_BIT_ALGN_MOVE_0_sqmuxa_2_i (.A(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_1_Z), .B(
        un1_restart_trng_fg_10_sn_1), .C(tap_cnt_0_sqmuxa_1_Z), .Y(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_i_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[71]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[71]), .C(
        un10_early_flags[71]), .Y(late_flags_7_fast_0[71]));
    SLE \no_early_no_late_val_end2[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[2]));
    SLE \late_flags[66]  (.D(late_flags_7_fast_0[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[66]));
    CFG4 #( .INIT(16'h1101) )  \bitalign_curr_state_34_4_0_.m37_0  (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[0]), .C(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .D(BIT_ALGN_ERR_c), .Y(m37));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_179  (.A(
        late_flags_Z[91]), .B(late_flags_Z[90]), .C(late_flags_Z[89]), 
        .D(late_flags_Z[88]), .Y(calc_done25_179));
    ARI1 #( .INIT(20'h48200) )  tapcnt_final_upd_8_s_6 (.A(VCC), .B(
        N_12_i), .C(tap_cnt_Z[6]), .D(tapcnt_final_upd_1_sqmuxa), .FCI(
        tapcnt_final_upd_8_cry_5), .S(tapcnt_final_upd_8[6]), .Y(
        tapcnt_final_upd_8_s_6_Y_0), .FCO(tapcnt_final_upd_8_s_6_FCO_0)
        );
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_12 (.A(
        early_flags_pmux_63_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[36]), .D(early_flags_Z[100]), .FCI(
        early_flags_pmux_63_1_1_co0_5), .S(
        early_flags_pmux_63_1_1_wmux_12_S_0), .Y(
        early_flags_pmux_63_1_1_y1_0), .FCO(
        early_flags_pmux_63_1_1_co1_5));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[4]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[4]), .C(
        un10_early_flags[4]), .Y(early_flags_7_fast_0[4]));
    SLE \tapcnt_final[3]  (.D(tapcnt_final_13_1_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[3]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_10 (.A(
        early_flags_pmux_126_1_0_0_y21), .B(
        early_flags_pmux_126_1_0_0_y9), .C(emflag_cnt_Z[2]), .D(VCC), 
        .FCI(early_flags_pmux_126_1_0_co0_4), .S(
        early_flags_pmux_126_1_0_wmux_10_S_0), .Y(
        early_flags_pmux_126_1_0_wmux_10_Y_0), .FCO(
        early_flags_pmux_126_1_0_co1_4));
    CFG2 #( .INIT(4'h8) )  bitalign_curr_state152_3 (.A(
        bitalign_curr_state152_1_Z), .B(bitalign_curr_state148_2_Z), 
        .Y(bitalign_curr_state152_3_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_27 (.A(
        un10_early_flags_2_0[24]), .B(un10_early_flags_1_Z[24]), .C(
        un10_early_flags_1_Z[3]), .Y(un10_early_flags[27]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_11 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[11]));
    CFG4 #( .INIT(16'hFFC8) )  un1_bitalign_curr_state_0_sqmuxa_9_4 (
        .A(calc_done28), .B(bitalign_curr_state162_Z), .C(calc_done27), 
        .D(un1_bitalign_curr_state_0_sqmuxa_9_2_Z), .Y(
        un1_bitalign_curr_state_0_sqmuxa_9_4_Z));
    SLE \bitalign_curr_state[3]  (.D(bitalign_curr_state_34[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[3]));
    SLE \tapcnt_final_upd[3]  (.D(tapcnt_final_upd_8[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[3]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_120 (.A(tap_cnt_Z[2]), 
        .B(un10_early_flags_1_Z[0]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[120]));
    SLE \late_flags[30]  (.D(late_flags_7_fast_0[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[30]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_73 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_Z[69]), .C(
        un10_early_flags_2_0[72]), .Y(un10_early_flags[73]));
    SLE \late_flags[51]  (.D(late_flags_7_fast_0[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[51]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[9]), 
        .D(early_flags_Z[73]), .FCI(early_flags_pmux_126_1_1_co1_0), 
        .S(early_flags_pmux_126_1_1_wmux_3_S_0), .Y(
        early_flags_pmux_126_1_1_y0_1), .FCO(
        early_flags_pmux_126_1_1_co0_1));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_0 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[53]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[53]), .C(
        un10_early_flags[53]), .Y(late_flags_7_fast_0[53]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_6 (.A(
        un10_tapcnt_final_6), .B(early_late_diff_Z[6]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_5_Z), .S(
        un1_early_late_diff_cry_6_S_0), .Y(
        un1_early_late_diff_cry_6_Y_0), .FCO(
        un1_early_late_diff_cry_6_Z));
    CFG2 #( .INIT(4'h1) )  rx_trng_done1_2_sqmuxa_0_398_i_a5 (.A(
        mv_dn_fg_Z), .B(mv_up_fg_Z), .Y(N_1416));
    CFG4 #( .INIT(16'h2000) )  tapcnt_final_3_sqmuxa (.A(
        bitalign_curr_state162_Z), .B(un1_calc_done25_5), .C(
        tapcnt_final27), .D(un1_early_late_diff_valid_Z), .Y(
        tapcnt_final_3_sqmuxa_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_6 (.A(
        late_flags_pmux_126_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[59]), .D(late_flags_Z[123]), .FCI(
        late_flags_pmux_126_1_0_co0_2), .S(
        late_flags_pmux_126_1_0_wmux_6_S_0), .Y(
        late_flags_pmux_126_1_0_0_y7), .FCO(
        late_flags_pmux_126_1_0_co1_2));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_36 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[32]), .C(
        un10_early_flags_1_Z[36]), .Y(un10_early_flags[36]));
    CFG2 #( .INIT(4'hE) )  \bitalign_curr_state_34_4_0_.un34lto7_3  (
        .A(un16_tapcnt_final_6), .B(un16_tapcnt_final_7), .Y(
        un34lto7_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[32]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[32]), .C(
        un10_early_flags[32]), .Y(late_flags_7_fast_0[32]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[0]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[0]), .D(GND), .FCI(
        emflag_cnt_cry_cy), .S(emflag_cnt_s[0]), .Y(
        emflag_cnt_cry_Y_1[0]), .FCO(emflag_cnt_cry_Z[0]));
    CFG2 #( .INIT(4'h8) )  \tapcnt_final_13_1[6]  (.A(
        tapcnt_final_13_Z[6]), .B(un1_tapcnt_final_0_sqmuxa_Z), .Y(
        tapcnt_final_13_1_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[20]), 
        .D(late_flags_Z[84]), .FCI(late_flags_pmux_63_1_1_co1_5), .S(
        late_flags_pmux_63_1_1_wmux_13_S_0), .Y(
        late_flags_pmux_63_1_1_y0_5), .FCO(
        late_flags_pmux_63_1_1_co0_6));
    SLE \early_flags[115]  (.D(early_flags_7_fast_0[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[115]));
    SLE \late_flags[117]  (.D(late_flags_7_fast_0[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[117]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[103]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[103]), .C(
        un10_early_flags[103]), .Y(early_flags_7_fast_0[103]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[15]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[15]), .C(
        un10_early_flags[15]), .Y(late_flags_7_fast_0[15]));
    SLE \tapcnt_final[4]  (.D(tapcnt_final_13_1_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[22]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[22]), .C(
        un10_early_flags[22]), .Y(late_flags_7_fast_0[22]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[19]), 
        .D(early_flags_Z[83]), .FCI(early_flags_pmux_126_1_0_0_co1), 
        .S(early_flags_pmux_126_1_0_wmux_1_S_0), .Y(
        early_flags_pmux_126_1_0_y0_0), .FCO(
        early_flags_pmux_126_1_0_co0_0));
    CFG4 #( .INIT(16'h00CE) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNI91ETE  (
        .A(m86_1), .B(m85_1), .C(bitalign_curr_state_Z[3]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[2]));
    SLE \no_early_no_late_val_st1[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[1]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_151  (.A(
        early_flags_Z[43]), .B(early_flags_Z[42]), .C(
        early_flags_Z[41]), .D(early_flags_Z[40]), .Y(calc_done25_151));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_20_1 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[20]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_116 (.A(tap_cnt_Z[3]), 
        .B(un10_early_flags_1_Z[20]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[116]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[79]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[79]), .C(
        un10_early_flags[79]), .Y(early_flags_7_fast_0[79]));
    CFG2 #( .INIT(4'h2) )  early_flags_1_sqmuxa (.A(
        bitalign_curr_state153_Z), .B(BIT_ALGN_OOR_0_c), .Y(
        early_flags_1_sqmuxa_Z));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_1 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[0]), .D(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[1]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_7 (.A(
        late_flags_pmux_63_1_1_y7), .B(late_flags_pmux_63_1_1_y5), .C(
        emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co1_2), .S(
        late_flags_pmux_63_1_1_wmux_7_S_0), .Y(
        late_flags_pmux_63_1_1_y0_3), .FCO(
        late_flags_pmux_63_1_1_co0_3));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_26 (.A(
        un10_early_flags_1_Z[10]), .B(un10_early_flags_2_0[24]), .C(
        un10_early_flags_1_Z[16]), .Y(un10_early_flags[26]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_10 (.A(
        un10_early_flags_1_Z[10]), .B(un10_early_flags_2_Z[10]), .C(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[10]));
    SLE \late_flags[61]  (.D(late_flags_7_fast_0[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[61]));
    SLE \early_flags[14]  (.D(early_flags_7_fast_0[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[14]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[91]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[91]), .C(
        un10_early_flags[91]), .Y(early_flags_7_fast_0[91]));
    CFG3 #( .INIT(8'hB1) )  \bitalign_curr_state_34_4_0_.m14  (.A(
        bitalign_curr_state_Z[2]), .B(N_8), .C(N_14), .Y(N_15));
    CFG4 #( .INIT(16'hFFFE) )  timeout_cnt_0_sqmuxa_RNIDBM31 (.A(
        restart_trng_fg_i), .B(timeout_cnt_0_sqmuxa_Z), .C(
        bitalign_curr_state_1_sqmuxa_7), .D(rx_err_1_sqmuxa_Z), .Y(
        timeout_cnte));
    ARI1 #( .INIT(20'h4AA00) )  rst_cnt_s_715 (.A(VCC), .B(
        rst_cnt_Z[0]), .C(GND), .D(GND), .FCI(VCC), .S(
        rst_cnt_s_715_S_0), .Y(rst_cnt_s_715_Y_0), .FCO(
        rst_cnt_s_715_FCO_0));
    SLE \no_early_no_late_val_st2[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[110]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[110]), .C(
        un10_early_flags[110]), .Y(late_flags_7_fast_0[110]));
    SLE \rst_cnt[3]  (.D(rst_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[73]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[73]), .C(
        un10_early_flags[73]), .Y(late_flags_7_fast_0[73]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[42]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[42]), .C(
        un10_early_flags[42]), .Y(late_flags_7_fast_0[42]));
    SLE \late_flags[25]  (.D(late_flags_7_fast_0[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[25]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[110]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[110]), .C(
        un10_early_flags[110]), .Y(early_flags_7_fast_0[110]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_2 (.A(
        un16_tapcnt_final_2), .B(early_late_diff_Z[2]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_1_Z), .S(
        un1_early_late_diff_1_cry_2_S_0), .Y(
        un1_early_late_diff_1_cry_2_Y_0), .FCO(
        un1_early_late_diff_1_cry_2_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[10]), 
        .D(late_flags_Z[74]), .FCI(late_flags_pmux_63_1_0_co1_0), .S(
        late_flags_pmux_63_1_0_wmux_3_S_0), .Y(
        late_flags_pmux_63_1_0_y0_1), .FCO(
        late_flags_pmux_63_1_0_co0_1));
    SLE \early_flags[49]  (.D(early_flags_RNO_0[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[49]));
    CFG4 #( .INIT(16'hFFFE) )  
        \bitalign_curr_state_34_4_0_.un2_noearly_nolate_diff_start_validlto7_2  
        (.A(un10_tapcnt_final_7), .B(un10_tapcnt_final_6), .C(
        un10_tapcnt_final_5), .D(un10_tapcnt_final_4), .Y(
        un2_noearly_nolate_diff_start_validlto7_2));
    CFG4 #( .INIT(16'h8000) )  rx_BIT_ALGN_ERR_4 (.A(timeout_cnt_Z[3]), 
        .B(timeout_cnt_Z[2]), .C(timeout_cnt_Z[1]), .D(
        timeout_cnt_Z[0]), .Y(rx_BIT_ALGN_ERR_4_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[7]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[7]), .C(
        un10_early_flags[7]), .Y(late_flags_7_fast_0[7]));
    ARI1 #( .INIT(20'h574B8) )  \tapcnt_final_RNIC3R56[5]  (.A(
        tap_cnt_Z[5]), .B(un1_tap_cnt_0_sqmuxa_14_0_0[1]), .C(N_60), 
        .D(tapcnt_final_Z[5]), .FCI(tap_cnt_17_i_m2_cry_4), .S(N_75), 
        .Y(tapcnt_final_RNIC3R56_Y_0[5]), .FCO(tap_cnt_17_i_m2_cry_5));
    CFG4 #( .INIT(16'h0800) )  
        \bitalign_curr_state_34_4_0_.calc_done25_253  (.A(
        calc_done25_236), .B(calc_done25_237), .C(calc_done25_253_1_0), 
        .D(calc_done25_245), .Y(calc_done25_253));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[4]  (.A(N_76), .B(N_63_0), .Y(
        N_24_i));
    SLE \noearly_nolate_diff_nxt[4]  (.D(noearly_nolate_diff_nxt_8[4]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_4));
    SLE \late_flags[106]  (.D(late_flags_7_fast_0[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[106]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_45 (.A(
        un10_early_flags_2_0[44]), .B(un10_early_flags_1_Z[40]), .C(
        un10_early_flags_1_Z[5]), .Y(un10_early_flags[45]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_106 (.A(
        un10_early_flags_1_Z[10]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[96]), .D(un10_early_flags_2_Z[10]), .Y(
        un10_early_flags[106]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[115]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[115]), .C(
        un10_early_flags[115]), .Y(late_flags_7_fast_0[115]));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_1_wmux_8 (.A(
        early_flags_pmux_126_1_1_y0_3), .B(early_flags_pmux_126_1_1_y3)
        , .C(early_flags_pmux_126_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_1_co0_3), .S(
        early_flags_pmux_126_1_1_wmux_8_S_0), .Y(
        early_flags_pmux_126_1_1_y9), .FCO(
        early_flags_pmux_126_1_1_co1_3));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_7 (.A(
        early_flags_pmux_126_1_0_0_y7), .B(
        early_flags_pmux_126_1_0_0_y5), .C(emflag_cnt_Z[4]), .D(
        emflag_cnt_Z[3]), .FCI(early_flags_pmux_126_1_0_co1_2), .S(
        early_flags_pmux_126_1_0_wmux_7_S_0), .Y(
        early_flags_pmux_126_1_0_y0_3), .FCO(
        early_flags_pmux_126_1_0_co0_3));
    SLE \early_flags[16]  (.D(early_flags_7_fast_0[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[16]));
    SLE \tapcnt_final[2]  (.D(tapcnt_final_13_1_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[2]));
    SLE \late_flags[87]  (.D(late_flags_7_fast_0[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[87]));
    SLE \early_flags[17]  (.D(early_flags_7_fast_0[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[17]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_180  (.A(
        late_flags_Z[79]), .B(late_flags_Z[78]), .C(late_flags_Z[77]), 
        .D(late_flags_Z[76]), .Y(calc_done25_180));
    CFG2 #( .INIT(4'hE) )  \tap_cnt_17_i_o2[6]  (.A(
        un1_bitalign_curr_state_1_sqmuxa_2_i_0), .B(restart_trng_fg_i), 
        .Y(N_63_0));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[107]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[107]), .C(
        un10_early_flags[107]), .Y(late_flags_7_fast_0[107]));
    SLE \early_flags[33]  (.D(early_flags_7_fast_0[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[33]));
    CFG4 #( .INIT(16'hECFE) )  un1_bitalign_curr_state_15_0 (.A(
        bitalign_curr_state_Z[1]), .B(un1_bitalign_curr_state_15_1_Z), 
        .C(bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state_15_0_Z));
    SLE late_last_set (.D(early_late_diff_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(late_last_set_Z));
    SLE \late_flags[75]  (.D(late_flags_7_fast_0[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[75]));
    CFG2 #( .INIT(4'h8) )  rx_BIT_ALGN_MOVE_0_sqmuxa_1 (.A(
        bitalign_curr_state156_Z), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_236  (.A(
        calc_done25_179), .B(calc_done25_178), .C(calc_done25_177), .D(
        calc_done25_176), .Y(calc_done25_236));
    SLE \early_flags[50]  (.D(early_flags_RNO_0[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[50]));
    CFG4 #( .INIT(16'h5504) )  \bitalign_curr_state_34_4_0_.m93  (.A(
        early_flags_dec[127]), .B(N_20), .C(late_last_set15_Z), .D(
        bitalign_curr_state_Z[0]), .Y(N_94));
    CFG2 #( .INIT(4'h1) )  
        \bitalign_curr_state148.bitalign_curr_state148_3_1  (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state163_2));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_0_wmux_20 (.A(
        early_flags_pmux_63_1_0_y0_8), .B(early_flags_pmux_63_1_0_y3_0)
        , .C(early_flags_pmux_63_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co0_9), .S(
        early_flags_pmux_63_1_0_wmux_20_S_0), .Y(
        early_flags_pmux_63_1_0_0_y21), .FCO(
        early_flags_pmux_63_1_0_co1_9));
    SLE \early_flags[11]  (.D(early_flags_7_fast_0[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[11]));
    CFG4 #( .INIT(16'hFFC8) )  un1_bitalign_curr_state_0_sqmuxa_9_2 (
        .A(calc_done25), .B(bitalign_curr_state162_Z), .C(calc_done26), 
        .D(un1_bitalign_curr_state_0_sqmuxa_9_1_Z), .Y(
        un1_bitalign_curr_state_0_sqmuxa_9_2_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_3 (.A(
        un16_tapcnt_final_3), .B(early_late_diff_Z[3]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_2_Z), .S(
        un1_early_late_diff_1_cry_3_S_0), .Y(
        un1_early_late_diff_1_cry_3_Y_0), .FCO(
        un1_early_late_diff_1_cry_3_Z));
    SLE \no_early_no_late_val_end1[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[1]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[24]), 
        .D(early_flags_Z[88]), .FCI(early_flags_pmux_63_1_1_co1_1), .S(
        early_flags_pmux_63_1_1_wmux_5_S_0), .Y(
        early_flags_pmux_63_1_1_y0_2), .FCO(
        early_flags_pmux_63_1_1_co0_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[30]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[30]), .C(
        un10_early_flags[30]), .Y(early_flags_7_fast_0[30]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[59]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[59]), .C(
        un10_early_flags[59]), .Y(late_flags_7_fast_0[59]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_4 (.A(
        un10_tapcnt_final_4), .B(un16_tapcnt_final_4), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_3_Z), .S(
        un10_tapcnt_final_cry_4_S_0), .Y(un10_tapcnt_final_cry_4_Y_0), 
        .FCO(un10_tapcnt_final_cry_4_Z));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_5 (.A(
        tapcnt_final_upd_Z[5]), .B(tapcnt_final_Z[5]), .C(tap_cnt_Z[5])
        , .D(N_1416), .Y(bitalign_curr_state61_5_Z));
    SLE \late_flags[17]  (.D(late_flags_7_fast_0[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[17]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_153  (.A(
        early_flags_Z[19]), .B(early_flags_Z[18]), .C(
        early_flags_Z[17]), .D(early_flags_Z[16]), .Y(calc_done25_153));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[17]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[17]), .C(
        un10_early_flags[17]), .Y(late_flags_7_fast_0[17]));
    SLE \tapcnt_final[0]  (.D(tapcnt_final_13_1_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[18]), 
        .D(early_flags_Z[82]), .FCI(early_flags_pmux_63_1_0_0_co1), .S(
        early_flags_pmux_63_1_0_wmux_1_S_0), .Y(
        early_flags_pmux_63_1_0_y0_0), .FCO(
        early_flags_pmux_63_1_0_co0_0));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_84 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[64]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[4]), .Y(
        un10_early_flags[84]));
    SLE \late_flags[35]  (.D(late_flags_7_fast_0[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[35]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_141  (.A(
        early_flags_Z[67]), .B(early_flags_Z[66]), .C(
        early_flags_Z[65]), .D(early_flags_Z[64]), .Y(calc_done25_141));
    SLE \early_flags[25]  (.D(early_flags_7_fast_0[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[25]));
    CFG4 #( .INIT(16'h1302) )  \bitalign_curr_state_34_4_0_.m39  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[4]), .C(
        i12_mux_0), .D(N_31), .Y(N_40));
    CFG4 #( .INIT(16'hF0CA) )  \bitalign_curr_state_34_4_0_.m74_1_0  (
        .A(N_9), .B(N_11), .C(rx_err_Z), .D(bitalign_curr_state_Z[1]), 
        .Y(m74_1_0_0));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_1_0 (.A(
        emflag_cnt_Z[1]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[1]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_0), .S(
        noearly_nolate_diff_nxt_8[1]), .Y(
        noearly_nolate_diff_nxt_8_cry_1_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_1));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIGUQVD[3]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNINKIR_0[3]), .B(
        early_val_RNI6FJ81_Z[3]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[3]), .FCI(tapcnt_final_13_m1_cry_2), .S(
        tapcnt_final_13_m1[3]), .Y(early_val_RNIGUQVD_Y[3]), .FCO(
        tapcnt_final_13_m1_cry_3));
    SLE \early_flags[63]  (.D(early_flags_7_fast_0[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[63]));
    SLE \rst_cnt[6]  (.D(rst_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[6]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_118 (.A(tap_cnt_Z[3]), 
        .B(un10_early_flags_1_Z[6]), .C(un10_early_flags_1_Z[64]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[118]));
    CFG2 #( .INIT(4'h4) )  \tapcnt_final_upd_8[0]  (.A(
        mv_dn_fg_0_sqmuxa_i_o2_0), .B(tap_cnt_Z[0]), .Y(
        tapcnt_final_upd_8_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[52]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[52]), .C(
        un10_early_flags[52]), .Y(early_flags_7_fast_0[52]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[31]), 
        .D(late_flags_Z[95]), .FCI(late_flags_pmux_126_1_0_co1_7), .S(
        late_flags_pmux_126_1_0_wmux_17_S_0), .Y(
        late_flags_pmux_126_1_0_y0_7), .FCO(
        late_flags_pmux_126_1_0_co0_8));
    SLE \late_flags[47]  (.D(late_flags_7_fast_0[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[47]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_4 (.A(
        un16_tapcnt_final_4), .B(early_late_diff_Z[4]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_3_Z), .S(
        un1_early_late_diff_1_cry_4_S_0), .Y(
        un1_early_late_diff_1_cry_4_Y_0), .FCO(
        un1_early_late_diff_1_cry_4_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_52 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[32]), .C(
        un10_early_flags_2_0[52]), .Y(un10_early_flags[52]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_10 (.A(
        late_flags_pmux_126_1_1_y21), .B(late_flags_pmux_126_1_1_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_126_1_1_co0_4), .S(
        late_flags_pmux_126_1_1_wmux_10_S_0), .Y(
        late_flags_pmux_126_1_1_wmux_10_Y_0), .FCO(
        late_flags_pmux_126_1_1_co1_4));
    SLE \emflag_cnt[4]  (.D(emflag_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[34]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[34]), .C(
        un10_early_flags[34]), .Y(late_flags_7_fast_0[34]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI6FJ81[3]  (.A(early_val_Z[3])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[3]), .Y(
        early_val_RNI6FJ81_Z[3]));
    CFG2 #( .INIT(4'h4) )  bitalign_curr_state153_1 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state153_1_Z));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state148_5 (.A(
        bitalign_curr_state162_Z), .B(un1_bitalign_curr_state148_5_4_Z)
        , .C(bitalign_curr_state164_Z), .Y(
        un1_bitalign_curr_state148_5_Z));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_230  (.A(
        calc_done25_155), .B(calc_done25_154), .C(calc_done25_153), .D(
        calc_done25_152), .Y(calc_done25_230));
    SLE \late_flags[1]  (.D(late_flags_7_fast_0[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[1]));
    CFG3 #( .INIT(8'hE4) )  \early_flags_RNO[50]  (.A(N_209), .B(
        EYE_MONITOR_EARLY_net_0_0), .C(early_flags_Z[50]), .Y(
        early_flags_RNO_0[50]));
    CFG4 #( .INIT(16'h4073) )  \bitalign_curr_state_34_4_0_.m7_1_0  (
        .A(BIT_ALGN_OOR_0_c), .B(bitalign_curr_state_Z[0]), .C(
        bitalign_curr_state41_Z), .D(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .Y(
        m7_1_1));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_14 (.A(
        late_flags_pmux_63_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[54]), .D(late_flags_Z[118]), .FCI(
        late_flags_pmux_63_1_0_co0_6), .S(
        late_flags_pmux_63_1_0_wmux_14_S_0), .Y(
        late_flags_pmux_63_1_0_y3_0), .FCO(
        late_flags_pmux_63_1_0_co1_6));
    CFG2 #( .INIT(4'hE) )  un1_sig_re_train (.A(rx_trng_done_Z), .B(
        rx_trng_done1_Z), .Y(un1_sig_re_train_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_1 (.A(
        un16_tapcnt_final_1), .B(early_late_diff_Z[1]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_0_Z), .S(
        un1_early_late_diff_1_cry_1_S_0), .Y(
        un1_early_late_diff_1_cry_1_Y_0), .FCO(
        un1_early_late_diff_1_cry_1_Z));
    SLE \early_flags[106]  (.D(early_flags_7_fast_0[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[106]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[24]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[24]), .C(
        un10_early_flags[24]), .Y(late_flags_7_fast_0[24]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_12 (.A(
        late_flags_pmux_63_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[36]), .D(late_flags_Z[100]), .FCI(
        late_flags_pmux_63_1_1_co0_5), .S(
        late_flags_pmux_63_1_1_wmux_12_S_0), .Y(
        late_flags_pmux_63_1_1_y1_0), .FCO(
        late_flags_pmux_63_1_1_co1_5));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_152  (.A(
        early_flags_Z[23]), .B(early_flags_Z[22]), .C(
        early_flags_Z[21]), .D(early_flags_Z[20]), .Y(calc_done25_152));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIROIR[5]  (.A(
        late_val_Z[5]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[5]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIROIR_0[5]));
    SLE \early_flags[52]  (.D(early_flags_7_fast_0[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[52]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_48 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_1_Z[48]), .C(
        un10_early_flags_2_0[48]), .Y(un10_early_flags[48]));
    CFG2 #( .INIT(4'h2) )  tap_cnt_0_sqmuxa_1_0 (.A(
        tap_cnt_0_sqmuxa_0_Z), .B(bitalign_curr_state_Z[1]), .Y(
        tap_cnt_0_sqmuxa_1_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[85]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[85]), .C(
        un10_early_flags[85]), .Y(late_flags_7_fast_0[85]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_4 (.A(
        early_flags_pmux_126_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[43]), .D(early_flags_Z[107]), .FCI(
        early_flags_pmux_126_1_0_co0_1), .S(
        early_flags_pmux_126_1_0_wmux_4_S_0), .Y(
        early_flags_pmux_126_1_0_0_y5), .FCO(
        early_flags_pmux_126_1_0_co1_1));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_62 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_1_Z[32]), .Y(
        un10_early_flags[62]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[56]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[56]), .C(
        un10_early_flags[56]), .Y(late_flags_7_fast_0[56]));
    CFG3 #( .INIT(8'h40) )  rx_err_2_sqmuxa_0_373_a2 (.A(
        restart_trng_fg_i), .B(early_flags_dec[127]), .C(
        bitalign_curr_state162_Z), .Y(N_1392));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[9]), .D(
        late_flags_Z[73]), .FCI(late_flags_pmux_126_1_1_co1_0), .S(
        late_flags_pmux_126_1_1_wmux_3_S_0), .Y(
        late_flags_pmux_126_1_1_y0_1), .FCO(
        late_flags_pmux_126_1_1_co0_1));
    CFG4 #( .INIT(16'h0F0E) )  emflag_cnt_1_sqmuxa_1 (.A(
        bitalign_curr_state160_Z), .B(bitalign_curr_state159), .C(
        early_flags_dec[127]), .D(bitalign_curr_state161_Z), .Y(
        emflag_cnt_1_sqmuxa_1_Z));
    CFG4 #( .INIT(16'h8000) )  timeout_cnt_0_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state154_Z), 
        .C(rx_err_Z), .D(calc_done_Z), .Y(timeout_cnt_0_sqmuxa_Z));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[2]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[2]), .D(GND), .FCI(
        emflag_cnt_cry_Z[1]), .S(emflag_cnt_s[2]), .Y(
        emflag_cnt_cry_Y_1[2]), .FCO(emflag_cnt_cry_Z[2]));
    SLE rx_BIT_ALGN_DIR (.D(un1_restart_trng_fg_6_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_BIT_ALGN_DIR_0_sqmuxa_2_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[34]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[34]), .C(
        un10_early_flags[34]), .Y(early_flags_7_fast_0[34]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[42]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[42]), .C(
        un10_early_flags[42]), .Y(early_flags_7_fast_0[42]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI8J6J1[2]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[2]), .D(GND), .FCI(
        timeout_cnt_cry[1]), .S(timeout_cnt_s[2]), .Y(
        timeout_cnt_RNI8J6J1_Y_0[2]), .FCO(timeout_cnt_cry[2]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_5_0 (
        .A(emflag_cnt_Z[5]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[5]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_4), .S(
        noearly_nolate_diff_start_7[5]), .Y(
        noearly_nolate_diff_start_7_cry_5_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[79]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[79]), .C(
        un10_early_flags[79]), .Y(late_flags_7_fast_0[79]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[23]), 
        .D(early_flags_Z[87]), .FCI(early_flags_pmux_126_1_0_co1_5), 
        .S(early_flags_pmux_126_1_0_wmux_13_S_0), .Y(
        early_flags_pmux_126_1_0_y0_5), .FCO(
        early_flags_pmux_126_1_0_co0_6));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNIIHTC3[6]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[6]), .D(GND), .FCI(
        timeout_cnt_cry[5]), .S(timeout_cnt_s[6]), .Y(
        timeout_cnt_RNIIHTC3_Y_0[6]), .FCO(timeout_cnt_cry[6]));
    CFG2 #( .INIT(4'h1) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_0 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .Y(
        tap_cnt_0_sqmuxa_2_0));
    CFG2 #( .INIT(4'h8) )  bitalign_curr_state149_1 (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state149_1_Z));
    CFG4 #( .INIT(16'hFFFE) )  
        \bitalign_curr_state_34_4_0_.late_cur_set_0_sqmuxa_i  (.A(
        un1_restart_trng_fg_10_sn_1), .B(tap_cnt_0_sqmuxa_1_Z), .C(
        early_last_set_1_sqmuxa_1_3_Z), .D(
        un1_bitalign_curr_state_2_sqmuxa), .Y(late_cur_set_0_sqmuxa_i));
    CFG2 #( .INIT(4'hE) )  tapcnt_final_13_m0s2 (.A(
        un1_restart_trng_fg_10_sn), .B(un1_bitalign_curr_state_12_Z), 
        .Y(tapcnt_final_13_m0s2_0));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_0 (.A(
        early_flags_pmux_126_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[33]), .D(early_flags_Z[97]), .FCI(
        early_flags_pmux_126_1_1_co0), .S(
        early_flags_pmux_126_1_1_wmux_0_S_0), .Y(
        early_flags_pmux_126_1_1_y1), .FCO(
        early_flags_pmux_126_1_1_co1));
    CFG2 #( .INIT(4'h4) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89  (.A(
        early_flags_pmux), .B(late_flags_pmux), .Y(
        bitalign_curr_state89));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_6_0 (.A(
        emflag_cnt_Z[6]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[6]), .D(GND), .FCI(early_late_diff_8_cry_5), .S(
        early_late_diff_8[6]), .Y(early_late_diff_8_cry_6_0_Y_0), .FCO(
        early_late_diff_8_cry_6));
    SLE \early_flags[73]  (.D(early_flags_7_fast_0[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[73]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_1 (.A(
        un10_tapcnt_final_1), .B(un16_tapcnt_final_1), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_0_Z), .S(
        un10_tapcnt_final_cry_1_S_0), .Y(un10_tapcnt_final_cry_1_Y_0), 
        .FCO(un10_tapcnt_final_cry_1_Z));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_108 (.A(tap_cnt_Z[4]), 
        .B(un10_early_flags_1_Z[12]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[108]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNICLJ81[5]  (.A(early_val_Z[5])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[5]), .Y(
        early_val_RNICLJ81_Z[5]));
    CFG2 #( .INIT(4'hD) )  early_late_diff_0_sqmuxa_RNIDTT8 (.A(
        early_late_diff_0_sqmuxa_1_0_Z), .B(early_late_diff_0_sqmuxa_Z)
        , .Y(early_late_diff_0_sqmuxa_1_i));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_16 (.A(
        late_flags_pmux_126_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[45]), .D(late_flags_Z[109]), .FCI(
        late_flags_pmux_126_1_1_co0_7), .S(
        late_flags_pmux_126_1_1_wmux_16_S_0), .Y(
        late_flags_pmux_126_1_1_y5_0), .FCO(
        late_flags_pmux_126_1_1_co1_7));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_0 (.A(
        late_flags_pmux_126_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[33]), .D(late_flags_Z[97]), .FCI(
        late_flags_pmux_126_1_1_co0), .S(
        late_flags_pmux_126_1_1_wmux_0_S_0), .Y(
        late_flags_pmux_126_1_1_y1), .FCO(late_flags_pmux_126_1_1_co1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[44]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[44]), .C(
        un10_early_flags[44]), .Y(late_flags_7_fast_0[44]));
    SLE \tap_cnt[5]  (.D(N_1497_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tap_cnt_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[127]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[127]), .C(
        un10_early_flags[127]), .Y(late_flags_7_fast_0[127]));
    CFG4 #( .INIT(16'h0BFB) )  \bitalign_curr_state_34_4_0_.m46  (.A(
        un1_retrain_adj_tap_i), .B(bitalign_curr_state13), .C(
        bitalign_curr_state_Z[0]), .D(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(N_47));
    CFG4 #( .INIT(16'h0010) )  rx_trng_done1_RNO (.A(restart_trng_fg_i)
        , .B(N_1416), .C(bitalign_curr_state_Z[3]), .D(
        bitalign_curr_state_Z[2]), .Y(N_1415_i));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[71]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[71]), .C(
        un10_early_flags[71]), .Y(early_flags_7_fast_0[71]));
    ARI1 #( .INIT(20'h5D872) )  
        \un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11[0]  (.A(tap_cnt_Z[0]), 
        .B(N_60), .C(N_89), .D(tapcnt_final_Z[0]), .FCI(GND), .S(
        un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_S_0[0]), .Y(
        un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_Y_0[0]), .FCO(
        tap_cnt_17_i_m2_cry_0));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_2_sqmuxa_1_0_a2 (.A(
        tapcnt_final_upd_1_sqmuxa), .B(restart_trng_fg_i), .Y(
        tapcnt_final_upd_2_sqmuxa_1));
    CFG3 #( .INIT(8'h51) )  \bitalign_curr_state_34_4_0_.m59  (.A(
        early_flags_dec[127]), .B(late_flags_pmux), .C(
        early_flags_pmux), .Y(N_60_0));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_229  (.A(
        calc_done25_151), .B(calc_done25_150), .C(calc_done25_149), .D(
        calc_done25_148), .Y(calc_done25_229));
    SLE \early_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_6 (.A(
        early_flags_pmux_126_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[57]), .D(early_flags_Z[121]), .FCI(
        early_flags_pmux_126_1_1_co0_2), .S(
        early_flags_pmux_126_1_1_wmux_6_S_0), .Y(
        early_flags_pmux_126_1_1_y7), .FCO(
        early_flags_pmux_126_1_1_co1_2));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_18 (.A(
        late_flags_pmux_126_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[63]), .D(late_flags_Z[127]), .FCI(
        late_flags_pmux_126_1_0_co0_8), .S(
        late_flags_pmux_126_1_0_wmux_18_S_0), .Y(
        late_flags_pmux_126_1_0_y7_0), .FCO(
        late_flags_pmux_126_1_0_co1_8));
    SLE \early_flags[80]  (.D(early_flags_7_fast_0[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[80]));
    CFG2 #( .INIT(4'h8) )  
        \bitalign_curr_state_34_4_0_.un2_noearly_nolate_diff_start_validlto1  
        (.A(un10_tapcnt_final_0), .B(un10_tapcnt_final_1), .Y(
        un2_noearly_nolate_diff_start_validlt2));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[25]), 
        .D(late_flags_Z[89]), .FCI(late_flags_pmux_126_1_1_co1_1), .S(
        late_flags_pmux_126_1_1_wmux_5_S_0), .Y(
        late_flags_pmux_126_1_1_y0_2), .FCO(
        late_flags_pmux_126_1_1_co0_2));
    SLE \late_flags[97]  (.D(late_flags_7_fast_0[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[97]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_3_0 (
        .A(emflag_cnt_Z[3]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[3]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_2), .S(
        noearly_nolate_diff_start_7[3]), .Y(
        noearly_nolate_diff_start_7_cry_3_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_3));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI99K12[3]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[3]), .D(GND), .FCI(
        timeout_cnt_cry[2]), .S(timeout_cnt_s[3]), .Y(
        timeout_cnt_RNI99K12_Y_0[3]), .FCO(timeout_cnt_cry[3]));
    CFG3 #( .INIT(8'hCD) )  calc_done_0_sqmuxa_2_i (.A(
        un1_bitalign_curr_state148_8_1_Z), .B(restart_trng_fg_i), .C(
        un1_bitalign_curr_state148_8_2_Z), .Y(calc_done_0_sqmuxa_2_i_Z)
        );
    SLE \noearly_nolate_diff_start[4]  (.D(
        noearly_nolate_diff_start_7[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_4));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_127_1_0_wmux (.A(
        emflag_cnt_Z[1]), .B(emflag_cnt_Z[0]), .C(
        late_flags_pmux_63_1_1_wmux_10_Y_0), .D(
        late_flags_pmux_63_1_0_wmux_10_Y_0), .FCI(VCC), .S(
        late_flags_pmux_127_1_0_wmux_S_0), .Y(
        late_flags_pmux_127_1_0_y0), .FCO(late_flags_pmux_127_1_0_co0));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_169  (.A(
        late_flags_Z[43]), .B(late_flags_Z[42]), .C(late_flags_Z[41]), 
        .D(late_flags_Z[40]), .Y(calc_done25_169));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_143  (.A(
        early_flags_Z[75]), .B(early_flags_Z[74]), .C(
        early_flags_Z[73]), .D(early_flags_Z[72]), .Y(calc_done25_143));
    CFG4 #( .INIT(16'h5150) )  sig_rx_BIT_ALGN_CLR_FLGS_11_iv (.A(
        restart_trng_fg_i), .B(rx_err_Z), .C(
        un1_bitalign_curr_state_1_sqmuxa_6_i_0), .D(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .Y(
        sig_rx_BIT_ALGN_CLR_FLGS_11));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNILLPT[1]  (.A(
        no_early_no_late_val_st1_Z[1]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[1]), .Y(
        un1_no_early_no_late_val_st1_1_1[1]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_18 (.A(
        early_flags_pmux_126_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[63]), .D(early_flags_Z[127]), .FCI(
        early_flags_pmux_126_1_0_co0_8), .S(
        early_flags_pmux_126_1_0_wmux_18_S_0), .Y(
        early_flags_pmux_126_1_0_y7_0), .FCO(
        early_flags_pmux_126_1_0_co1_8));
    SLE \early_flags[112]  (.D(early_flags_7_fast_0[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[112]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_12 (.A(
        late_flags_pmux_126_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[37]), .D(late_flags_Z[101]), .FCI(
        late_flags_pmux_126_1_1_co0_5), .S(
        late_flags_pmux_126_1_1_wmux_12_S_0), .Y(
        late_flags_pmux_126_1_1_y1_0), .FCO(
        late_flags_pmux_126_1_1_co1_5));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[4]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[4]), .D(GND), .FCI(
        emflag_cnt_cry_Z[3]), .S(emflag_cnt_s[4]), .Y(
        emflag_cnt_cry_Y_1[4]), .FCO(emflag_cnt_cry_Z[4]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[8]), 
        .D(early_flags_Z[72]), .FCI(early_flags_pmux_63_1_1_co1_0), .S(
        early_flags_pmux_63_1_1_wmux_3_S_0), .Y(
        early_flags_pmux_63_1_1_y0_1), .FCO(
        early_flags_pmux_63_1_1_co0_1));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_14 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[3]), .C(un10_early_flags_1_Z[6]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[14]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_185  (.A(
        late_flags_Z[115]), .B(late_flags_Z[114]), .C(
        late_flags_Z[113]), .D(late_flags_Z[112]), .Y(calc_done25_185));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_41 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_0[40]), .C(
        un10_early_flags_2_Z[37]), .Y(un10_early_flags[41]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[5]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[5]), .D(GND), .FCI(
        emflag_cnt_cry_Z[4]), .S(emflag_cnt_s[5]), .Y(
        emflag_cnt_cry_Y_1[5]), .FCO(emflag_cnt_cry_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[76]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[76]), .C(
        un10_early_flags[76]), .Y(late_flags_7_fast_0[76]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_16 (.A(
        late_flags_pmux_63_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[44]), .D(late_flags_Z[108]), .FCI(
        late_flags_pmux_63_1_1_co0_7), .S(
        late_flags_pmux_63_1_1_wmux_16_S_0), .Y(
        late_flags_pmux_63_1_1_y5_0), .FCO(
        late_flags_pmux_63_1_1_co1_7));
    SLE \late_flags[58]  (.D(late_flags_7_fast_0[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[58]));
    SLE \late_flags[108]  (.D(late_flags_7_fast_0[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[108]));
    CFG3 #( .INIT(8'hDC) )  un1_early_flags_1_sqmuxa_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(early_flags_1_sqmuxa_Z), .C(
        bitalign_curr_state156_Z), .Y(un1_early_flags_1_sqmuxa_1_Z));
    SLE \early_flags[18]  (.D(early_flags_7_fast_0[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[18]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[111]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[111]), .C(
        un10_early_flags[111]), .Y(late_flags_7_fast_0[111]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_188  (.A(
        late_flags_Z[103]), .B(late_flags_Z[102]), .C(
        late_flags_Z[101]), .D(late_flags_Z[100]), .Y(calc_done25_188));
    SLE \rst_cnt[1]  (.D(rst_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[1]));
    CFG3 #( .INIT(8'h20) )  bitalign_curr_state_1_sqmuxa_7_0_a2 (.A(
        un1_retrain_adj_tap_i), .B(bitalign_curr_state12_Z), .C(N_98), 
        .Y(bitalign_curr_state_1_sqmuxa_7));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_110 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[64]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_1_Z[40]), .Y(
        un10_early_flags[110]));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state148_5_4 (.A(
        bitalign_curr_state154_3_Z), .B(bitalign_curr_state149_Z), .C(
        bitalign_curr_state148_Z), .Y(un1_bitalign_curr_state148_5_4_Z)
        );
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_10 (.A(
        early_flags_pmux_63_1_1_y21), .B(early_flags_pmux_63_1_1_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_63_1_1_co0_4), .S(
        early_flags_pmux_63_1_1_wmux_10_S_0), .Y(
        early_flags_pmux_63_1_1_wmux_10_Y_0), .FCO(
        early_flags_pmux_63_1_1_co1_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[100]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[100]), .C(
        un10_early_flags[100]), .Y(early_flags_7_fast_0[100]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_55 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_47_0_Z), .Y(
        un10_early_flags[55]));
    SLE \early_flags[90]  (.D(early_flags_7_fast_0[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[90]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_142  (.A(
        early_flags_Z[79]), .B(early_flags_Z[78]), .C(
        early_flags_Z[77]), .D(early_flags_Z[76]), .Y(calc_done25_142));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_1_wmux_8 (.A(
        late_flags_pmux_63_1_1_y0_3), .B(late_flags_pmux_63_1_1_y3), 
        .C(late_flags_pmux_63_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co0_3), .S(
        late_flags_pmux_63_1_1_wmux_8_S_0), .Y(
        late_flags_pmux_63_1_1_y9), .FCO(late_flags_pmux_63_1_1_co1_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[10]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[10]), .C(
        un10_early_flags[10]), .Y(late_flags_7_fast_0[10]));
    ARI1 #( .INIT(20'h400DC) )  \emflag_cnt_cry_cy[0]  (.A(
        un1_restart_trng_fg_9_0_443_0), .B(bitalign_curr_state_Z[0]), 
        .C(bitalign_curr_state_Z[2]), .D(bitalign_curr_state_Z[4]), 
        .FCI(VCC), .S(emflag_cnt_cry_cy_S_1[0]), .Y(
        emflag_cnt_cry_cy_Y_1[0]), .FCO(emflag_cnt_cry_cy));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[87]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[87]), .C(
        un10_early_flags[87]), .Y(late_flags_7_fast_0[87]));
    SLE \late_flags[83]  (.D(late_flags_7_fast_0[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[83]));
    SLE \early_flags[82]  (.D(early_flags_7_fast_0[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[82]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_87 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_3_Z[87]), .Y(
        un10_early_flags[87]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_139  (.A(
        early_flags_Z[91]), .B(early_flags_Z[90]), .C(
        early_flags_Z[89]), .D(early_flags_Z[88]), .Y(calc_done25_139));
    CFG2 #( .INIT(4'h2) )  
        \bitalign_curr_state_34_4_0_.late_cur_set_2_sqmuxa  (.A(
        un1_bitalign_curr_state_2_sqmuxa), .B(restart_trng_fg_i), .Y(
        late_cur_set_2_sqmuxa));
    SLE \wait_cnt[0]  (.D(wait_cnt_4_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(wait_cnt_Z[0]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_0 (.A(
        un16_tapcnt_final_0), .B(un10_tapcnt_final_0), .C(GND), .D(GND)
        , .FCI(GND), .S(un16_tapcnt_final_cry_0_S_0), .Y(
        un16_tapcnt_final_cry_0_Y_0), .FCO(un16_tapcnt_final_cry_0_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[57]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[57]), .C(
        un10_early_flags[57]), .Y(early_flags_7_fast_0[57]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_4 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_2_0[0]), .D(
        un10_early_flags_2_Z[4]), .Y(un10_early_flags[4]));
    SLE \no_early_no_late_val_st1[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[6]));
    SLE \late_flags[68]  (.D(late_flags_7_fast_0[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[68]));
    CFG2 #( .INIT(4'h1) )  \bitalign_curr_state_34_4_0_.m8  (.A(
        bitalign_curr_state_Z[0]), .B(BIT_ALGN_OOR_0_c), .Y(N_9));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_65 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[6]), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[65]));
    CFG3 #( .INIT(8'h80) )  early_late_diff_0_sqmuxa (.A(
        late_flags_pmux), .B(late_last_set15_Z), .C(
        bitalign_curr_state161_Z), .Y(early_late_diff_0_sqmuxa_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_40 (.A(
        un10_early_flags_2_0[40]), .B(un10_early_flags_1_Z[0]), .C(
        un10_early_flags_1_Z[40]), .Y(un10_early_flags[40]));
    CFG4 #( .INIT(16'hFFFE) )  early_last_set_0_sqmuxa_i (.A(
        un1_restart_trng_fg_10_sn_1), .B(early_last_set_1_sqmuxa_1_3_Z)
        , .C(early_val_0_sqmuxa_1_0_Z), .D(tap_cnt_0_sqmuxa_1_Z), .Y(
        early_last_set_0_sqmuxa_i_Z));
    SLE \early_late_diff[4]  (.D(early_late_diff_8[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[4]));
    CFG4 #( .INIT(16'hFFCE) )  un1_bitalign_curr_state_16_1 (.A(
        bitalign_curr_state_Z[2]), .B(un1_bitalign_curr_state_14_1_Z), 
        .C(bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[4]), .Y(
        un1_bitalign_curr_state_16_1_Z));
    SLE \late_flags[13]  (.D(late_flags_7_fast_0[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[13]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_126_1_0_co1_3), .S(
        late_flags_pmux_126_1_0_wmux_9_S_0), .Y(
        late_flags_pmux_126_1_0_wmux_9_Y_0), .FCO(
        late_flags_pmux_126_1_0_co0_4));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[95]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[95]), .C(
        un10_early_flags[95]), .Y(late_flags_7_fast_0[95]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_47_0 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[6]), .Y(un10_early_flags_47_0_Z));
    SLE \timeout_cnt[6]  (.D(timeout_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[6]));
    SLE \tap_cnt[1]  (.D(N_30_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[1]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_2 (.A(
        late_flags_pmux_63_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[50]), .D(late_flags_Z[114]), .FCI(
        late_flags_pmux_63_1_0_co0_0), .S(
        late_flags_pmux_63_1_0_wmux_2_S_0), .Y(
        late_flags_pmux_63_1_0_0_y3), .FCO(
        late_flags_pmux_63_1_0_co1_0));
    CFG3 #( .INIT(8'h20) )  \bitalign_curr_state_34_4_0_.m66_2  (.A(
        bitalign_curr_state_Z[3]), .B(bitalign_curr_state_Z[4]), .C(
        N_65), .Y(m66_1));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[6]  (.A(
        no_early_no_late_val_end1_Z[6]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[6]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[20]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[20]), .C(
        un10_early_flags[20]), .Y(early_flags_7_fast_0[20]));
    SLE \early_flags[3]  (.D(early_flags_7_fast_0[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[3]));
    CFG4 #( .INIT(16'hFF9C) )  \wait_cnt_4[1]  (.A(wait_cnt_Z[0]), .B(
        wait_cnt_Z[1]), .C(bitalign_curr_state152_3_Z), .D(
        un1_restart_trng_fg_0), .Y(wait_cnt_4_Z[1]));
    CFG2 #( .INIT(4'hD) )  early_val_0_sqmuxa_1_i (.A(
        early_cur_set_0_sqmuxa_1_Z), .B(un1_tap_cnt_0_sqmuxa_6_0), .Y(
        early_val_0_sqmuxa_1_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[80]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[80]), .C(
        un10_early_flags[80]), .Y(early_flags_7_fast_0[80]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_100 (.A(
        un10_early_flags_1_Z[36]), .B(un10_early_flags_1_Z[64]), .C(
        un10_early_flags_2_0[100]), .Y(un10_early_flags[100]));
    CFG2 #( .INIT(4'h8) )  sig_rx_BIT_ALGN_CLR_FLGS14 (.A(CO0_0), .B(
        cnt_Z[1]), .Y(sig_rx_BIT_ALGN_CLR_FLGS14_Z));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_0_0 (.A(
        emflag_cnt_Z[0]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[0]), .D(GND), .FCI(early_late_diff_8_cry_0_0_cy_Z), 
        .S(early_late_diff_8[0]), .Y(early_late_diff_8_cry_0_0_Y_0), 
        .FCO(early_late_diff_8_cry_0));
    CFG4 #( .INIT(16'h8000) )  early_flags_dec_127 (.A(emflag_cnt_Z[2])
        , .B(early_flags_dec_127_4_Z), .C(emflag_cnt_Z[1]), .D(
        emflag_cnt_Z[0]), .Y(early_flags_dec[127]));
    SLE \late_flags[54]  (.D(late_flags_7_fast_0[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[54]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_2 (.A(
        early_flags_pmux_126_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[49]), .D(early_flags_Z[113]), .FCI(
        early_flags_pmux_126_1_1_co0_0), .S(
        early_flags_pmux_126_1_1_wmux_2_S_0), .Y(
        early_flags_pmux_126_1_1_y3), .FCO(
        early_flags_pmux_126_1_1_co1_0));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_170  (.A(
        late_flags_Z[39]), .B(late_flags_Z[38]), .C(late_flags_Z[37]), 
        .D(late_flags_Z[36]), .Y(calc_done25_170));
    SLE \late_flags[43]  (.D(late_flags_7_fast_0[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[43]));
    SLE \early_flags[92]  (.D(early_flags_7_fast_0[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[92]));
    CFG3 #( .INIT(8'h08) )  bitalign_curr_state_1_sqmuxa_4 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state149_Z), 
        .C(BIT_ALGN_ERR_c), .Y(bitalign_curr_state_1_sqmuxa_4_Z));
    SLE \early_flags[124]  (.D(early_flags_7_fast_0[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[124]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[47]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[47]), .C(
        un10_early_flags[47]), .Y(early_flags_7_fast_0[47]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_0_wmux_20 (.A(
        late_flags_pmux_63_1_0_y0_8), .B(late_flags_pmux_63_1_0_y3_0), 
        .C(late_flags_pmux_63_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co0_9), .S(
        late_flags_pmux_63_1_0_wmux_20_S_0), .Y(
        late_flags_pmux_63_1_0_0_y21), .FCO(
        late_flags_pmux_63_1_0_co1_9));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[15]), 
        .D(late_flags_Z[79]), .FCI(late_flags_pmux_126_1_0_co1_6), .S(
        late_flags_pmux_126_1_0_wmux_15_S_0), .Y(
        late_flags_pmux_126_1_0_y0_6), .FCO(
        late_flags_pmux_126_1_0_co0_7));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[60]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[60]), .C(
        un10_early_flags[60]), .Y(early_flags_7_fast_0[60]));
    CFG2 #( .INIT(4'h6) )  \cnt_RNO[1]  (.A(CO0_0), .B(cnt_Z[1]), .Y(
        cnt_RNO_0[1]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_86 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[6]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[6]), .Y(
        un10_early_flags[86]));
    SLE \early_flags[45]  (.D(early_flags_7_fast_0[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[45]));
    CFG4 #( .INIT(16'hAE00) )  
        \bitalign_curr_state_34_4_0_.tapcnt_final_2_sqmuxa  (.A(
        calc_done28), .B(calc_done27), .C(un10_tapcnt_final_cry_7_Z), 
        .D(bitalign_curr_state162_Z), .Y(tapcnt_final_2_sqmuxa));
    CFG3 #( .INIT(8'h46) )  \bitalign_curr_state_34_4_0_.m12  (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state_Z[0]), 
        .C(bitalign_curr_state61), .Y(N_114_mux));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_100_2_0 (.A(
        un10_early_flags_2_Z[4]), .B(tap_cnt_Z[4]), .Y(
        un10_early_flags_2_0[100]));
    SLE \late_flags[122]  (.D(late_flags_7_fast_0[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[122]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_16_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[3]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[16]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_58 (.A(tap_cnt_Z[6]), 
        .B(un10_early_flags_1_Z[10]), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[58]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[62]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[62]), .C(
        un10_early_flags[62]), .Y(late_flags_7_fast_0[62]));
    CFG4 #( .INIT(16'hFFBA) )  un1_bitalign_curr_state_15_2 (.A(
        un1_bitalign_curr_state_15_0_Z), .B(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .C(bitalign_curr_state155), .D(
        early_flags_0_sqmuxa_Z), .Y(un1_bitalign_curr_state_15_2_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_18 (.A(
        late_flags_pmux_63_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[62]), .D(late_flags_Z[126]), .FCI(
        late_flags_pmux_63_1_0_co0_8), .S(
        late_flags_pmux_63_1_0_wmux_18_S_0), .Y(
        late_flags_pmux_63_1_0_y7_0), .FCO(
        late_flags_pmux_63_1_0_co1_8));
    CFG3 #( .INIT(8'hB1) )  \bitalign_curr_state_34_4_0_.m13  (.A(
        bitalign_curr_state_Z[1]), .B(N_11), .C(N_114_mux), .Y(N_14));
    CFG4 #( .INIT(16'h0040) )  bitalign_curr_state164 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state152_1_Z), .D(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state164_Z));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[1]  (.A(N_79), .B(N_63_0), .Y(
        N_30_i));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_24_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[2]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[24]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_19 (.A(
        early_flags_pmux_63_1_1_y7_0), .B(early_flags_pmux_63_1_1_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co1_8), .S(
        early_flags_pmux_63_1_1_wmux_19_S_0), .Y(
        early_flags_pmux_63_1_1_y0_8), .FCO(
        early_flags_pmux_63_1_1_co0_9));
    SLE \late_flags[22]  (.D(late_flags_7_fast_0[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[22]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_7 (.A(
        un16_tapcnt_final_7), .B(un10_tapcnt_final_7), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_6_Z), .S(
        un16_tapcnt_final_cry_7_S_0), .Y(un16_tapcnt_final_cry_7_Y_0), 
        .FCO(un16_tapcnt_final_cry_7_Z));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[2]  (.A(
        no_early_no_late_val_end1_Z[2]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[2]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[2]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_3 (.A(
        un10_tapcnt_final_3), .B(un16_tapcnt_final_3), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_2_Z), .S(
        un10_tapcnt_final_cry_3_S_0), .Y(un10_tapcnt_final_cry_3_Y_0), 
        .FCO(un10_tapcnt_final_cry_3_Z));
    CFG4 #( .INIT(16'h0400) )  un10_early_flags_79 (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[6]), .C(tap_cnt_Z[5]), .D(
        un10_early_flags_1_0[15]), .Y(un10_early_flags[79]));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.m43_0_a2_0  (
        .A(BIT_ALGN_ERR_c), .B(retrain_reg_Z[2]), .Y(
        un1_rx_BIT_ALGN_START));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[1]  (.A(
        no_early_no_late_val_end1_Z[1]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[1]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[1]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_4 (.A(
        late_flags_pmux_126_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[43]), .D(late_flags_Z[107]), .FCI(
        late_flags_pmux_126_1_0_co0_1), .S(
        late_flags_pmux_126_1_0_wmux_4_S_0), .Y(
        late_flags_pmux_126_1_0_0_y5), .FCO(
        late_flags_pmux_126_1_0_co1_1));
    CFG4 #( .INIT(16'h72AA) )  \bitalign_curr_state_34_4_0_.m30  (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state41_Z), .C(
        bit_align_dly_done_Z), .D(bitalign_curr_state_Z[1]), .Y(N_31));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[23]), 
        .D(late_flags_Z[87]), .FCI(late_flags_pmux_126_1_0_co1_5), .S(
        late_flags_pmux_126_1_0_wmux_13_S_0), .Y(
        late_flags_pmux_126_1_0_y0_5), .FCO(
        late_flags_pmux_126_1_0_co0_6));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_68 (.A(tap_cnt_Z[2]), 
        .B(tap_cnt_Z[6]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[68]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_14 (.A(
        late_flags_pmux_63_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[52]), .D(late_flags_Z[116]), .FCI(
        late_flags_pmux_63_1_1_co0_6), .S(
        late_flags_pmux_63_1_1_wmux_14_S_0), .Y(
        late_flags_pmux_63_1_1_y3_0), .FCO(
        late_flags_pmux_63_1_1_co1_6));
    SLE \late_flags[64]  (.D(late_flags_7_fast_0[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[64]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[7]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[7]), .C(
        un10_early_flags[7]), .Y(early_flags_7_fast_0[7]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[24]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[24]), .C(
        un10_early_flags[24]), .Y(early_flags_7_fast_0[24]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[84]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[84]), .C(
        un10_early_flags[84]), .Y(early_flags_7_fast_0[84]));
    SLE \no_early_no_late_val_st1[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[59]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[59]), .C(
        un10_early_flags[59]), .Y(early_flags_7_fast_0[59]));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_3_sqmuxa_1_0_a2 (.A(
        tapcnt_final_upd_2_sqmuxa), .B(restart_trng_fg_i), .Y(
        tapcnt_final_upd_3_sqmuxa_1));
    CFG4 #( .INIT(16'hFFF8) )  un1_bitalign_curr_state_1_sqmuxa_2 (.A(
        tap_cnt_0_sqmuxa_1_0_Z), .B(tap_cnt_0_sqmuxa_2_0), .C(
        bitalign_curr_state_1_sqmuxa_4_Z), .D(tap_cnt_0_sqmuxa_1_Z), 
        .Y(un1_bitalign_curr_state_1_sqmuxa_2_i_0));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNITTPT[5]  (.A(
        no_early_no_late_val_st1_Z[5]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[5]), .Y(
        un1_no_early_no_late_val_st1_1_1[5]));
    CFG3 #( .INIT(8'h40) )  un10_early_flags_17 (.A(N_1498), .B(
        un10_early_flags_2_Z[8]), .C(un10_early_flags_2_0[16]), .Y(
        un10_early_flags[17]));
    SLE \late_flags[72]  (.D(late_flags_7_fast_0[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[72]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_0 (.A(
        early_flags_pmux_63_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[32]), .D(early_flags_Z[96]), .FCI(
        early_flags_pmux_63_1_1_co0), .S(
        early_flags_pmux_63_1_1_wmux_0_S_0), .Y(
        early_flags_pmux_63_1_1_y1), .FCO(early_flags_pmux_63_1_1_co1));
    SLE \timeout_cnt[0]  (.D(timeout_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[0]));
    SLE \late_flags[114]  (.D(late_flags_7_fast_0[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[114]));
    SLE \late_flags[3]  (.D(late_flags_7_fast_0[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[3]));
    SLE \late_flags[100]  (.D(late_flags_7_fast_0[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[100]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[18]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[18]), .C(
        un10_early_flags[18]), .Y(late_flags_7_fast_0[18]));
    CFG4 #( .INIT(16'hDDEC) )  \bitalign_curr_state_34_4_0_.m91  (.A(
        bitalign_curr_state_Z[2]), .B(m91_1), .C(N_116_mux), .D(
        m91_1_0), .Y(N_92));
    CFG4 #( .INIT(16'hFEFC) )  mv_dn_fg_0_sqmuxa_i_o2 (.A(
        bitalign_curr_state148_Z), .B(bitalign_curr_state_1_sqmuxa_4_Z)
        , .C(restart_trng_fg_i), .D(N_61), .Y(mv_dn_fg_0_sqmuxa_i_o2_0)
        );
    CFG4 #( .INIT(16'hFDFC) )  un1_restart_trng_fg_8 (.A(
        early_flags_pmux), .B(un1_tap_cnt_0_sqmuxa_6_0), .C(
        restart_trng_fg_i), .D(early_val_0_sqmuxa_1_0_Z), .Y(
        un1_restart_trng_fg_8_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[64]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[64]), .C(
        un10_early_flags[64]), .Y(early_flags_7_fast_0[64]));
    SLE \late_flags[93]  (.D(late_flags_7_fast_0[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[93]));
    SLE \late_flags[89]  (.D(late_flags_7_fast_0[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[89]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[38]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[38]), .C(
        un10_early_flags[38]), .Y(early_flags_7_fast_0[38]));
    ARI1 #( .INIT(20'h574B8) )  \tapcnt_final_RNISU155[4]  (.A(
        tap_cnt_Z[4]), .B(un1_tap_cnt_0_sqmuxa_14_0_0[1]), .C(N_60), 
        .D(tapcnt_final_Z[4]), .FCI(tap_cnt_17_i_m2_cry_3), .S(N_76), 
        .Y(tapcnt_final_RNISU155_Y_0[4]), .FCO(tap_cnt_17_i_m2_cry_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[123]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[123]), .C(
        un10_early_flags[123]), .Y(early_flags_7_fast_0[123]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_32_2_0 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[32]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[97]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[97]), .C(
        un10_early_flags[97]), .Y(late_flags_7_fast_0[97]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_51 (.A(
        un10_early_flags_1_Z[3]), .B(un10_early_flags_2_0[48]), .C(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[51]));
    SLE \late_flags[32]  (.D(late_flags_7_fast_0[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[32]));
    CFG2 #( .INIT(4'hE) )  un1_bitalign_curr_state_15_1 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[4]), .Y(
        un1_bitalign_curr_state_15_1_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[8]  (.A(VCC), .B(
        rst_cnt_Z[8]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[7]), .S(
        rst_cnt_s[8]), .Y(rst_cnt_cry_Y_1[8]), .FCO(rst_cnt_cry_Z[8]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_7 (.A(
        late_flags_pmux_63_1_0_0_y7), .B(late_flags_pmux_63_1_0_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co1_2), .S(
        late_flags_pmux_63_1_0_wmux_7_S_0), .Y(
        late_flags_pmux_63_1_0_y0_3), .FCO(
        late_flags_pmux_63_1_0_co0_3));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[16]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[16]), .C(
        un10_early_flags[16]), .Y(early_flags_7_fast_0[16]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[35]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[35]), .C(
        un10_early_flags[35]), .Y(early_flags_7_fast_0[35]));
    CFG3 #( .INIT(8'h1B) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNIAODV4  (
        .A(bitalign_curr_state_Z[0]), .B(m82_1_0), .C(m82_1_1), .Y(
        N_83));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_10_2 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[10]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_0 (.A(late_val_Z[0])
        , .B(early_val_Z[0]), .C(GND), .D(GND), .FCI(GND), .S(
        tapcnt_final27_cry_0_S_0), .Y(tapcnt_final27_cry_0_Y_0), .FCO(
        tapcnt_final27_cry_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[80]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[80]), .C(
        un10_early_flags[80]), .Y(late_flags_7_fast_0[80]));
    SLE \late_flags[119]  (.D(late_flags_7_fast_0[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[119]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_67_2 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[67]));
    CFG4 #( .INIT(16'h8000) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(tap_cnt_0_sqmuxa_2_0), .C(
        bitalign_curr_state_Z[1]), .D(un1_bitalign_curr_state151_Z), 
        .Y(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_Z));
    SLE \late_flags[9]  (.D(late_flags_7_fast_0[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[9]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[5]  (.A(
        tapcnt_final_Z[5]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[5]), .Y(
        tapcnt_final_13_Z[5]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIJTRFA[2]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNILIIR_0[2]), .B(
        early_val_RNI3CJ81_Z[2]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[2]), .FCI(tapcnt_final_13_m1_cry_1), .S(
        tapcnt_final_13_m1[2]), .Y(early_val_RNIJTRFA_Y[2]), .FCO(
        tapcnt_final_13_m1_cry_2));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[6]), 
        .D(early_flags_Z[70]), .FCI(early_flags_pmux_63_1_0_co1_4), .S(
        early_flags_pmux_63_1_0_wmux_11_S_0), .Y(
        early_flags_pmux_63_1_0_y0_4), .FCO(
        early_flags_pmux_63_1_0_co0_5));
    SLE \late_flags[19]  (.D(late_flags_7_fast_0[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[19]));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_6 (.A(
        tapcnt_final_upd_Z[6]), .B(tapcnt_final_Z[6]), .C(tap_cnt_Z[6])
        , .D(N_1416), .Y(bitalign_curr_state61_6_Z));
    CFG4 #( .INIT(16'h0800) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state_2_sqmuxa_4_0  
        (.A(bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), 
        .C(early_flags_dec[127]), .D(
        bitalign_curr_state_2_sqmuxa_4_0_0), .Y(emflag_cnt_0_sqmuxa));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[3]  (.A(
        no_early_no_late_val_end1_Z[3]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[3]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[3]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIS2TV6[1]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIJGIR_0[1]), .B(
        early_val_RNI09J81_Z[1]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[1]), .FCI(tapcnt_final_13_m1_cry_0), .S(
        tapcnt_final_13_m1[1]), .Y(early_val_RNIS2TV6_Y[1]), .FCO(
        tapcnt_final_13_m1_cry_1));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_72_2_0 (.A(tap_cnt_Z[2]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[5]), .Y(
        un10_early_flags_2_0[72]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_61 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_2_Z[37]), .Y(
        un10_early_flags[61]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_19 (.A(
        late_flags_pmux_126_1_1_y7_0), .B(late_flags_pmux_126_1_1_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co1_8), .S(
        late_flags_pmux_126_1_1_wmux_19_S_0), .Y(
        late_flags_pmux_126_1_1_y0_8), .FCO(
        late_flags_pmux_126_1_1_co0_9));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[28]), 
        .D(late_flags_Z[92]), .FCI(late_flags_pmux_63_1_1_co1_7), .S(
        late_flags_pmux_63_1_1_wmux_17_S_0), .Y(
        late_flags_pmux_63_1_1_y0_7), .FCO(
        late_flags_pmux_63_1_1_co0_8));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_16 (.A(
        un10_early_flags_1_Z[16]), .B(un10_early_flags_2_Z[8]), .C(
        un10_early_flags_2_0[16]), .Y(un10_early_flags[16]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_231  (.A(
        calc_done25_159), .B(calc_done25_158), .C(calc_done25_157), .D(
        calc_done25_156), .Y(calc_done25_231));
    CFG4 #( .INIT(16'h1F0E) )  \bitalign_curr_state_34_4_0_.m50  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        m50_1_1), .D(N_47), .Y(N_51));
    SLE \early_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[1]));
    CFG4 #( .INIT(16'hFFFE) )  un2_noearly_nolate_diff_nxt_validlto7_2 
        (.A(un16_tapcnt_final_7), .B(un16_tapcnt_final_6), .C(
        un16_tapcnt_final_5), .D(un16_tapcnt_final_4), .Y(
        un2_noearly_nolate_diff_nxt_validlto7_2_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[2]  (.A(VCC), .B(
        rst_cnt_Z[2]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[1]), .S(
        rst_cnt_s[2]), .Y(rst_cnt_cry_Y_1[2]), .FCO(rst_cnt_cry_Z[2]));
    SLE \early_flags[24]  (.D(early_flags_7_fast_0[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[24]));
    SLE \late_flags[49]  (.D(late_flags_RNO_0[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[49]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[13]), 
        .D(late_flags_Z[77]), .FCI(late_flags_pmux_126_1_1_co1_6), .S(
        late_flags_pmux_126_1_1_wmux_15_S_0), .Y(
        late_flags_pmux_126_1_1_y0_6), .FCO(
        late_flags_pmux_126_1_1_co0_7));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_124 (.A(
        un10_early_flags_1_Z[12]), .B(tap_cnt_Z[1]), .C(
        un10_early_flags_1_Z[48]), .D(un10_early_flags_1_Z[64]), .Y(
        un10_early_flags[124]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_225  (.A(
        calc_done25_135), .B(calc_done25_134), .C(calc_done25_133), .D(
        calc_done25_132), .Y(calc_done25_225));
    CFG3 #( .INIT(8'hE0) )  \wait_cnt_4_RNO[2]  (.A(wait_cnt_Z[1]), .B(
        wait_cnt_Z[0]), .C(bitalign_curr_state152_3_Z), .Y(CO1));
    CFG4 #( .INIT(16'h0001) )  bitalign_curr_state61_0_0_RNIQOA01 (.A(
        bitalign_curr_state61_0), .B(bitalign_curr_state61_NE_4_Z), .C(
        bitalign_curr_state61_5_Z), .D(bitalign_curr_state61_4_Z), .Y(
        bitalign_curr_state61));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_4_2 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[4]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_127_1_0_wmux_0 (.A(
        early_flags_pmux_127_1_0_y0), .B(emflag_cnt_Z[0]), .C(
        early_flags_pmux_126_1_1_wmux_10_Y_0), .D(
        early_flags_pmux_126_1_0_wmux_10_Y_0), .FCI(
        early_flags_pmux_127_1_0_co0), .S(
        early_flags_pmux_127_1_0_wmux_0_S_0), .Y(early_flags_pmux), 
        .FCO(early_flags_pmux_127_1_0_co1));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_175  (.A(
        late_flags_Z[51]), .B(late_flags_Z[50]), .C(late_flags_Z[49]), 
        .D(late_flags_Z[48]), .Y(calc_done25_175));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_5 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_2_Z[4]), .Y(un10_early_flags[5]));
    SLE \early_flags[116]  (.D(early_flags_7_fast_0[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[116]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[8]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[8]), .C(
        un10_early_flags[8]), .Y(early_flags_7_fast_0[8]));
    CFG3 #( .INIT(8'h1D) )  \tapcnt_final_13_RNO_1[6]  (.A(
        no_early_no_late_val_st1_Z[6]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[6]), .Y(
        un1_no_early_no_late_val_st1_1_1[6]));
    SLE \no_early_no_late_val_st2[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[6]));
    CFG4 #( .INIT(16'hEDDE) )  \wait_cnt_4[2]  (.A(wait_cnt_Z[2]), .B(
        un1_restart_trng_fg_0), .C(bitalign_curr_state152_3_Z), .D(CO1)
        , .Y(wait_cnt_4_Z[2]));
    ARI1 #( .INIT(20'h54411) )  tapcnt_final_upd_8_cry_4_0 (.A(
        tap_cnt_Z[4]), .B(mv_dn_fg_0_sqmuxa_i_o2_0), .C(
        tapcnt_final_upd_1_sqmuxa), .D(GND), .FCI(
        tapcnt_final_upd_8_cry_3), .S(tapcnt_final_upd_8[4]), .Y(
        tapcnt_final_upd_8_cry_4_0_Y_0), .FCO(tapcnt_final_upd_8_cry_4)
        );
    CFG4 #( .INIT(16'hFFF6) )  un1_bitalign_curr_state_14_1_0 (.A(
        bitalign_curr_state_Z[3]), .B(bitalign_curr_state_Z[2]), .C(
        un1_bitalign_curr_state_14_1_Z), .D(
        tapcnt_final_upd_3_sqmuxa_Z), .Y(
        un1_bitalign_curr_state_14_1_0_Z));
    SLE \emflag_cnt[5]  (.D(emflag_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[5]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_178  (.A(
        late_flags_Z[95]), .B(late_flags_Z[94]), .C(late_flags_Z[93]), 
        .D(late_flags_Z[92]), .Y(calc_done25_178));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_0_wmux_8 (.A(
        late_flags_pmux_126_1_0_y0_3), .B(late_flags_pmux_126_1_0_0_y3)
        , .C(late_flags_pmux_126_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co0_3), .S(
        late_flags_pmux_126_1_0_wmux_8_S_0), .Y(
        late_flags_pmux_126_1_0_0_y9), .FCO(
        late_flags_pmux_126_1_0_co1_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[64]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[64]), .C(
        un10_early_flags[64]), .Y(late_flags_7_fast_0[64]));
    CFG3 #( .INIT(8'hCD) )  \bitalign_curr_state_34_4_0_.m37  (.A(
        m37_1_1), .B(m37), .C(early_flags_dec[127]), .Y(i12_mux_0));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_44 (.A(
        un10_early_flags_2_0[44]), .B(un10_early_flags_1_Z[32]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[44]));
    SLE \early_flags[13]  (.D(early_flags_7_fast_0[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[13]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_6 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_2_Z[6]), .Y(un10_early_flags[6]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNINNPT[2]  (.A(
        no_early_no_late_val_st1_Z[2]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[2]), .Y(
        un1_no_early_no_late_val_st1_1_1[2]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[14]), 
        .D(late_flags_Z[78]), .FCI(late_flags_pmux_63_1_0_co1_6), .S(
        late_flags_pmux_63_1_0_wmux_15_S_0), .Y(
        late_flags_pmux_63_1_0_y0_6), .FCO(
        late_flags_pmux_63_1_0_co0_7));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[90]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[90]), .C(
        un10_early_flags[90]), .Y(early_flags_7_fast_0[90]));
    CFG4 #( .INIT(16'hA0A3) )  \bitalign_curr_state_34_4_0_.m7  (.A(
        m7_1_1), .B(bitalign_curr_state12_Z), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        N_8));
    SLE \tap_cnt[4]  (.D(N_24_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[4]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIJJPT[0]  (.A(
        no_early_no_late_val_st1_Z[0]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[0]), .Y(
        un1_no_early_no_late_val_st1_1_1[0]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_60 (.A(tap_cnt_Z[6]), 
        .B(un10_early_flags_1_Z[12]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[60]));
    SLE \early_flags[26]  (.D(early_flags_7_fast_0[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[26]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_93 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[69]), .Y(
        un10_early_flags[93]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_10_1 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_1_Z[10]));
    SLE \early_flags[27]  (.D(early_flags_7_fast_0[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[27]));
    CFG4 #( .INIT(16'h0015) )  early_cur_set_0_sqmuxa_1 (.A(
        restart_trng_fg_i), .B(un1_early_last_set_1_sqmuxa_1_1_tz_Z), 
        .C(early_flags_pmux), .D(early_last_set_1_sqmuxa_1_3_Z), .Y(
        early_cur_set_0_sqmuxa_1_Z));
    SLE \late_flags[115]  (.D(late_flags_7_fast_0[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[115]));
    CFG2 #( .INIT(4'h4) )  \tapcnt_final_upd_8[1]  (.A(
        mv_dn_fg_0_sqmuxa_i_o2_0), .B(tap_cnt_Z[1]), .Y(
        tapcnt_final_upd_8_Z[1]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_52_2_0 (.A(
        un10_early_flags_2_Z[4]), .B(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[52]));
    SLE \tap_cnt[3]  (.D(N_26_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[3]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[19]), 
        .D(late_flags_Z[83]), .FCI(late_flags_pmux_126_1_0_0_co1), .S(
        late_flags_pmux_126_1_0_wmux_1_S_0), .Y(
        late_flags_pmux_126_1_0_y0_0), .FCO(
        late_flags_pmux_126_1_0_co0_0));
    SLE \early_flags[59]  (.D(early_flags_7_fast_0[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[59]));
    CFG2 #( .INIT(4'h1) )  bitalign_curr_state161_2 (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state161_2_Z));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_69_2 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[69]));
    SLE \timeout_cnt[2]  (.D(timeout_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[2]));
    SLE \no_early_no_late_val_end1[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[5]));
    CFG2 #( .INIT(4'h2) )  early_flags_1_sqmuxa_1 (.A(
        bitalign_curr_state148_Z), .B(bitalign_curr_state12_Z), .Y(
        early_flags_1_sqmuxa_1_Z));
    SLE \early_flags[21]  (.D(early_flags_7_fast_0[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[21]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[1]  (.A(
        tapcnt_final_Z[1]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[1]), .Y(
        tapcnt_final_13_Z[1]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_159  (.A(
        early_flags_Z[3]), .B(early_flags_Z[2]), .C(early_flags_Z[1]), 
        .D(early_flags_Z[0]), .Y(calc_done25_159));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_nxt_8_cry_0_0_cy (
        .A(VCC), .B(un1_restart_trng_fg_5_0), .C(GND), .D(GND), .FCI(
        VCC), .S(noearly_nolate_diff_nxt_8_cry_0_0_cy_S_0), .Y(
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_19 (.A(
        early_flags_pmux_63_1_0_y7_0), .B(early_flags_pmux_63_1_0_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co1_8), .S(
        early_flags_pmux_63_1_0_wmux_19_S_0), .Y(
        early_flags_pmux_63_1_0_y0_8), .FCO(
        early_flags_pmux_63_1_0_co0_9));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[3]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[3]), .C(
        un10_early_flags[3]), .Y(late_flags_7_fast_0[3]));
    SLE early_cur_set (.D(early_val_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_cur_set_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(early_cur_set_Z));
    SLE \retrain_reg[1]  (.D(retrain_reg_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(retrain_reg_Z[1]));
    CFG4 #( .INIT(16'h0020) )  bitalign_curr_state161 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state161_2_Z), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state161_Z));
    SLE \late_flags[99]  (.D(late_flags_7_fast_0[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[99]));
    CFG3 #( .INIT(8'h04) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNI46NMB  (
        .A(un1_bitalign_curr_state_0_sqmuxa_9_i), .B(N_102), .C(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[3]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[6]  (.A(
        tapcnt_final_Z[6]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[6]), .Y(
        tapcnt_final_13_Z[6]));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_0_0 (.A(
        tapcnt_final_upd_Z[0]), .B(tapcnt_final_Z[0]), .C(tap_cnt_Z[0])
        , .D(N_1416), .Y(bitalign_curr_state61_0));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[88]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[88]), .C(
        un10_early_flags[88]), .Y(late_flags_7_fast_0[88]));
    SLE \rst_cnt[8]  (.D(rst_cnt_s[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[8]));
    CFG4 #( .INIT(16'h0053) )  \bitalign_curr_state_34_4_0_.m49  (.A(
        N_9), .B(N_11), .C(rx_err_Z), .D(bitalign_curr_state_Z[1]), .Y(
        N_50));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[4]), .D(
        late_flags_Z[68]), .FCI(late_flags_pmux_63_1_1_co1_4), .S(
        late_flags_pmux_63_1_1_wmux_11_S_0), .Y(
        late_flags_pmux_63_1_1_y0_4), .FCO(
        late_flags_pmux_63_1_1_co0_5));
    SLE \late_flags[103]  (.D(late_flags_7_fast_0[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[103]));
    CFG3 #( .INIT(8'h40) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNIAJUD  (
        .A(early_flags_dec[127]), .B(bitalign_curr_state89), .C(
        bitalign_curr_state_Z[0]), .Y(N_108));
    CFG4 #( .INIT(16'h0010) )  bitalign_curr_state148 (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state148_2_Z), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state148_Z));
    CFG3 #( .INIT(8'hF6) )  \wait_cnt_4[0]  (.A(
        bitalign_curr_state152_3_Z), .B(wait_cnt_Z[0]), .C(
        un1_restart_trng_fg_0), .Y(wait_cnt_4_Z[0]));
    CFG2 #( .INIT(4'hD) )  bit_align_done_0_sqmuxa_3_i (.A(
        bit_align_done_0_sqmuxa_3_1_Z), .B(bit_align_done_0_sqmuxa_2_Z)
        , .Y(bit_align_done_0_sqmuxa_3_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[33]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[33]), .C(
        un10_early_flags[33]), .Y(early_flags_7_fast_0[33]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[3]  (.A(
        tapcnt_final_Z[3]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[3]), .Y(
        tapcnt_final_13_Z[3]));
    CFG4 #( .INIT(16'hEA00) )  
        \bitalign_curr_state_34_4_0_.tapcnt_final_1_sqmuxa_2  (.A(
        calc_done26), .B(calc_done27), .C(un10_tapcnt_final_cry_7_Z), 
        .D(bitalign_curr_state162_Z), .Y(tapcnt_final_1_sqmuxa_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[51]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[51]), .C(
        un10_early_flags[51]), .Y(early_flags_7_fast_0[51]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[16]), 
        .D(early_flags_Z[80]), .FCI(early_flags_pmux_63_1_1_co1), .S(
        early_flags_pmux_63_1_1_wmux_1_S_0), .Y(
        early_flags_pmux_63_1_1_y0_0), .FCO(
        early_flags_pmux_63_1_1_co0_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[94]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[94]), .C(
        un10_early_flags[94]), .Y(early_flags_7_fast_0[94]));
    CFG4 #( .INIT(16'h3332) )  bit_align_start_RNO (.A(sig_re_train_Z), 
        .B(restart_trng_fg_i), .C(bit_align_done_0_sqmuxa_2_Z), .D(
        bitalign_curr_state_1_sqmuxa_4_Z), .Y(N_1439_i));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[90]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[90]), .C(
        un10_early_flags[90]), .Y(late_flags_7_fast_0[90]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[35]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[35]), .C(
        un10_early_flags[35]), .Y(late_flags_7_fast_0[35]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_122 (.A(tap_cnt_Z[2]), 
        .B(un10_early_flags_1_Z[10]), .C(un10_early_flags_1_Z[64]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[122]));
    CFG4 #( .INIT(16'h2772) )  \tapcnt_final_13_RNO_0[6]  (.A(
        tapcnt_final_3_sqmuxa_Z), .B(late_val_Z[6]), .C(
        un1_no_early_no_late_val_end1_1_1_Z[6]), .D(
        un1_no_early_no_late_val_st1_1_1[6]), .Y(
        tapcnt_final_13_m1_axb_6_1));
    SLE \early_flags[107]  (.D(early_flags_7_fast_0[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[107]));
    CFG4 #( .INIT(16'hFFFE) )  
        \bitalign_curr_state_34_4_0_.un34lto7_4  (.A(
        un16_tapcnt_final_3), .B(un16_tapcnt_final_2), .C(
        un16_tapcnt_final_1), .D(un16_tapcnt_final_0), .Y(un34lto7_4));
    CFG4 #( .INIT(16'h8000) )  reset_dly_fg4 (.A(rst_cnt_Z[0]), .B(
        reset_dly_fg4_8_Z), .C(rst_cnt_Z[1]), .D(reset_dly_fg4_4_Z), 
        .Y(reset_dly_fg4_Z));
    SLE \late_flags[101]  (.D(late_flags_7_fast_0[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[101]));
    CFG1 #( .INIT(2'h1) )  tapcnt_final_upd_8_s_6_RNO (.A(
        mv_dn_fg_0_sqmuxa_i_o2_0), .Y(N_12_i));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[25]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[25]), .C(
        un10_early_flags[25]), .Y(late_flags_7_fast_0[25]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_3_0 (.A(
        emflag_cnt_Z[3]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[3]), .D(GND), .FCI(early_late_diff_8_cry_2), .S(
        early_late_diff_8[3]), .Y(early_late_diff_8_cry_3_0_Y_0), .FCO(
        early_late_diff_8_cry_3));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[2]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[2]), .C(
        un10_early_flags[2]), .Y(early_flags_7_fast_0[2]));
    SLE \early_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[2]));
    CFG4 #( .INIT(16'hCCEC) )  mv_dn_fg_0_sqmuxa_i_0 (.A(N_98), .B(
        mv_dn_fg_0_sqmuxa_i_o2_0), .C(mv_up_fg_Z), .D(mv_dn_fg_Z), .Y(
        mv_dn_fg_0_sqmuxa_i_0_0));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_160  (.A(
        late_flags_Z[15]), .B(late_flags_Z[14]), .C(late_flags_Z[13]), 
        .D(late_flags_Z[12]), .Y(calc_done25_160));
    SLE \no_early_no_late_val_st2[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[4]));
    SLE \tap_cnt[2]  (.D(N_28_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[2]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_64_2_0 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[5]), .Y(
        un10_early_flags_2_0[64]));
    SLE bit_align_done (.D(bit_align_done_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        bit_align_done_0_sqmuxa_3_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(bit_align_done_Z)
        );
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[4]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[4]), .C(
        un10_early_flags[4]), .Y(late_flags_7_fast_0[4]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[3]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[3]), .C(
        un10_early_flags[3]), .Y(early_flags_7_fast_0[3]));
    CFG3 #( .INIT(8'h73) )  no_early_no_late_val_st1_0_sqmuxa_i (.A(
        un1_early_flags_pmux_1_Z), .B(early_late_diff_0_sqmuxa_1_0_Z), 
        .C(emflag_cnt_0_sqmuxa), .Y(
        no_early_no_late_val_st1_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[41]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[41]), .C(
        un10_early_flags[41]), .Y(early_flags_7_fast_0[41]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[102]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[102]), .C(
        un10_early_flags[102]), .Y(late_flags_7_fast_0[102]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[11]), 
        .D(early_flags_Z[75]), .FCI(early_flags_pmux_126_1_0_co1_0), 
        .S(early_flags_pmux_126_1_0_wmux_3_S_0), .Y(
        early_flags_pmux_126_1_0_y0_1), .FCO(
        early_flags_pmux_126_1_0_co0_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[28]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[28]), .C(
        un10_early_flags[28]), .Y(early_flags_7_fast_0[28]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[6]), .D(
        late_flags_Z[70]), .FCI(late_flags_pmux_63_1_0_co1_4), .S(
        late_flags_pmux_63_1_0_wmux_11_S_0), .Y(
        late_flags_pmux_63_1_0_y0_4), .FCO(
        late_flags_pmux_63_1_0_co0_5));
    CFG3 #( .INIT(8'hD0) )  early_flags_0_sqmuxa_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(BIT_ALGN_ERR_c), .C(
        bitalign_curr_state149_Z), .Y(early_flags_0_sqmuxa_1_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[88]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[88]), .C(
        un10_early_flags[88]), .Y(early_flags_7_fast_0[88]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_0_wmux_20 (.A(
        late_flags_pmux_126_1_0_y0_8), .B(late_flags_pmux_126_1_0_y3_0)
        , .C(late_flags_pmux_126_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co0_9), .S(
        late_flags_pmux_126_1_0_wmux_20_S_0), .Y(
        late_flags_pmux_126_1_0_0_y21), .FCO(
        late_flags_pmux_126_1_0_co1_9));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state148_4_1 (.A(
        bitalign_curr_state164_Z), .B(bitalign_curr_state162_Z), .C(
        bitalign_curr_state163_Z), .Y(un1_bitalign_curr_state148_4_1_Z)
        );
    CFG3 #( .INIT(8'hCE) )  mv_up_fg_0_sqmuxa_i_0 (.A(N_98), .B(
        mv_dn_fg_0_sqmuxa_i_o2_0), .C(mv_up_fg_Z), .Y(
        mv_up_fg_0_sqmuxa_i_0_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[25]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[25]), .C(
        un10_early_flags[25]), .Y(early_flags_7_fast_0[25]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[45]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[45]), .C(
        un10_early_flags[45]), .Y(late_flags_7_fast_0[45]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[2]  (.A(
        tapcnt_final_Z[2]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[2]), .Y(
        tapcnt_final_13_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[85]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[85]), .C(
        un10_early_flags[85]), .Y(early_flags_7_fast_0[85]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[30]), 
        .D(early_flags_Z[94]), .FCI(early_flags_pmux_63_1_0_co1_7), .S(
        early_flags_pmux_63_1_0_wmux_17_S_0), .Y(
        early_flags_pmux_63_1_0_y0_7), .FCO(
        early_flags_pmux_63_1_0_co0_8));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_0_wmux_8 (.A(
        early_flags_pmux_63_1_0_y0_3), .B(early_flags_pmux_63_1_0_0_y3)
        , .C(early_flags_pmux_63_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co0_3), .S(
        early_flags_pmux_63_1_0_wmux_8_S_0), .Y(
        early_flags_pmux_63_1_0_0_y9), .FCO(
        early_flags_pmux_63_1_0_co1_3));
    CFG3 #( .INIT(8'h20) )  bitalign_curr_state160 (.A(
        bitalign_curr_state152_1_Z), .B(bitalign_curr_state_Z[4]), .C(
        bitalign_curr_state149_1_Z), .Y(bitalign_curr_state160_Z));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_5 (.A(
        un10_tapcnt_final_5), .B(un16_tapcnt_final_5), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_4_Z), .S(
        un10_tapcnt_final_cry_5_S_0), .Y(un10_tapcnt_final_cry_5_Y_0), 
        .FCO(un10_tapcnt_final_cry_5_Z));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_6_2 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_2_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[68]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[68]), .C(
        un10_early_flags[68]), .Y(early_flags_7_fast_0[68]));
    SLE \early_flags[89]  (.D(early_flags_7_fast_0[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[89]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_149  (.A(
        early_flags_Z[35]), .B(early_flags_Z[34]), .C(
        early_flags_Z[33]), .D(early_flags_Z[32]), .Y(calc_done25_149));
    CFG2 #( .INIT(4'h1) )  \bitalign_curr_state_34_4_0_.m75  (.A(
        N_119_mux), .B(bitalign_curr_state_Z[0]), .Y(N_76_0));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_191  (.A(
        late_flags_Z[107]), .B(late_flags_Z[106]), .C(
        late_flags_Z[105]), .D(late_flags_Z[104]), .Y(calc_done25_191));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_6 (.A(
        un16_tapcnt_final_6), .B(un10_tapcnt_final_6), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_5_Z), .S(
        un16_tapcnt_final_cry_6_S_0), .Y(un16_tapcnt_final_cry_6_Y_0), 
        .FCO(un16_tapcnt_final_cry_6_Z));
    CFG4 #( .INIT(16'hFFF8) )  un1_early_last_set_1_sqmuxa_1_1_tz (.A(
        bitalign_curr_state160_Z), .B(early_cur_set_Z), .C(
        emflag_cnt_0_sqmuxa), .D(bitalign_curr_state159), .Y(
        un1_early_last_set_1_sqmuxa_1_1_tz_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[3]), .D(
        late_flags_Z[67]), .FCI(VCC), .S(
        late_flags_pmux_126_1_0_wmux_S_0), .Y(
        late_flags_pmux_126_1_0_0_y0), .FCO(
        late_flags_pmux_126_1_0_0_co0));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_2_0 (.A(
        emflag_cnt_Z[2]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[2]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_1), .S(
        noearly_nolate_diff_nxt_8[2]), .Y(
        noearly_nolate_diff_nxt_8_cry_2_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_2));
    SLE \noearly_nolate_diff_start[1]  (.D(
        noearly_nolate_diff_start_7[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_1));
    SLE \late_flags[50]  (.D(late_flags_RNO_0[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[50]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_130  (.A(
        early_flags_Z[127]), .B(early_flags_Z[126]), .C(
        early_flags_Z[125]), .D(early_flags_Z[124]), .Y(
        calc_done25_130));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[65]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[65]), .C(
        un10_early_flags[65]), .Y(early_flags_7_fast_0[65]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_47 (.A(
        un10_early_flags_47_0_Z), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[47]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[52]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[52]), .C(
        un10_early_flags[52]), .Y(late_flags_7_fast_0[52]));
    CFG4 #( .INIT(16'h8000) )  early_flags_dec_127_4 (.A(
        emflag_cnt_Z[4]), .B(emflag_cnt_Z[3]), .C(emflag_cnt_Z[6]), .D(
        emflag_cnt_Z[5]), .Y(early_flags_dec_127_4_Z));
    CFG4 #( .INIT(16'h8000) )  reset_dly_fg4_8 (.A(rst_cnt_Z[8]), .B(
        rst_cnt_Z[7]), .C(rst_cnt_Z[6]), .D(reset_dly_fg4_6_Z), .Y(
        reset_dly_fg4_8_Z));
    CFG3 #( .INIT(8'hEC) )  rx_trng_done1_1_sqmuxa_i_o2 (.A(
        un1_rx_BIT_ALGN_START), .B(bitalign_curr_state12_Z), .C(
        un1_retrain_adj_tap_i), .Y(N_61));
    CFG2 #( .INIT(4'h7) )  \bitalign_curr_state_34_4_0_.N_29_i  (.A(
        bitalign_curr_state41_Z), .B(bitalign_curr_state_Z[0]), .Y(
        N_29_i));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_33 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_2_0[32]), .Y(un10_early_flags[33]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[120]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[120]), .C(
        un10_early_flags[120]), .Y(early_flags_7_fast_0[120]));
    SLE \late_flags[126]  (.D(late_flags_7_fast_0[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[126]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[70]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[70]), .C(
        un10_early_flags[70]), .Y(early_flags_7_fast_0[70]));
    SLE \early_flags[28]  (.D(early_flags_7_fast_0[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[28]));
    SLE \restart_edge_reg[1]  (.D(restart_edge_reg_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[1]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_0_wmux_8 (.A(
        late_flags_pmux_63_1_0_y0_3), .B(late_flags_pmux_63_1_0_0_y3), 
        .C(late_flags_pmux_63_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co0_3), .S(
        late_flags_pmux_63_1_0_wmux_8_S_0), .Y(
        late_flags_pmux_63_1_0_0_y9), .FCO(
        late_flags_pmux_63_1_0_co1_3));
    SLE \early_late_diff[7]  (.D(early_late_diff_8[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[7]));
    SLE \no_early_no_late_val_st1[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[5]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_238  (.A(
        calc_done25_187), .B(calc_done25_186), .C(calc_done25_185), .D(
        calc_done25_184), .Y(calc_done25_238));
    SLE \early_flags[44]  (.D(early_flags_7_fast_0[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[44]));
    SLE \early_flags[121]  (.D(early_flags_7_fast_0[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[121]));
    CFG3 #( .INIT(8'hE4) )  \late_flags_RNO[50]  (.A(N_209), .B(
        EYE_MONITOR_LATE_net_0_0), .C(late_flags_Z[50]), .Y(
        late_flags_RNO_0[50]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[29]), 
        .D(early_flags_Z[93]), .FCI(early_flags_pmux_126_1_1_co1_7), 
        .S(early_flags_pmux_126_1_1_wmux_17_S_0), .Y(
        early_flags_pmux_126_1_1_y0_7), .FCO(
        early_flags_pmux_126_1_1_co0_8));
    CFG2 #( .INIT(4'h4) )  
        \bitalign_curr_state_34_4_0_.rx_BIT_ALGN_CLR_FLGS  (.A(
        rx_trng_done_Z), .B(sig_rx_BIT_ALGN_CLR_FLGS_Z), .Y(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_127_1_0_wmux_0 (.A(
        late_flags_pmux_127_1_0_y0), .B(emflag_cnt_Z[0]), .C(
        late_flags_pmux_126_1_1_wmux_10_Y_0), .D(
        late_flags_pmux_126_1_0_wmux_10_Y_0), .FCI(
        late_flags_pmux_127_1_0_co0), .S(
        late_flags_pmux_127_1_0_wmux_0_S_0), .Y(late_flags_pmux), .FCO(
        late_flags_pmux_127_1_0_co1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[37]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[37]), .C(
        un10_early_flags[37]), .Y(late_flags_7_fast_0[37]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_54 (.A(tap_cnt_Z[6]), 
        .B(un10_early_flags_2_Z[6]), .C(un10_early_flags_1_Z[6]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[54]));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[2]  (.A(N_78), .B(N_63_0), .Y(
        N_28_i));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_7 (.A(
        un10_tapcnt_final_7), .B(early_late_diff_Z[7]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_6_Z), .S(
        un1_early_late_diff_cry_7_S_0), .Y(
        un1_early_late_diff_cry_7_Y_0), .FCO(
        un1_early_late_diff_cry_7_Z));
    CFG3 #( .INIT(8'hFD) )  \tap_cnt_17_i_o2_0[6]  (.A(
        bitalign_curr_state_0_sqmuxa_10), .B(
        un1_early_flags_1_sqmuxa_i), .C(rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), 
        .Y(N_60));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[22]), 
        .D(late_flags_Z[86]), .FCI(late_flags_pmux_63_1_0_co1_5), .S(
        late_flags_pmux_63_1_0_wmux_13_S_0), .Y(
        late_flags_pmux_63_1_0_y0_5), .FCO(
        late_flags_pmux_63_1_0_co0_6));
    SLE \early_flags[99]  (.D(early_flags_7_fast_0[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[99]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_186  (.A(
        late_flags_Z[127]), .B(late_flags_Z[126]), .C(
        late_flags_Z[125]), .D(late_flags_Z[124]), .Y(calc_done25_186));
    CFG2 #( .INIT(4'h2) )  rx_trng_done_1_sqmuxa (.A(
        bitalign_curr_state164_Z), .B(bitalign_curr_state41_Z), .Y(
        rx_trng_done_1_sqmuxa_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[1]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[1]), .C(
        un10_early_flags[1]), .Y(early_flags_7_fast_0[1]));
    SLE \early_flags[100]  (.D(early_flags_7_fast_0[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[100]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_0 (.A(
        un16_tapcnt_final_0), .B(early_late_diff_Z[0]), .C(GND), .D(
        GND), .FCI(GND), .S(un1_early_late_diff_1_cry_0_S_0), .Y(
        un1_early_late_diff_1_cry_0_Y_0), .FCO(
        un1_early_late_diff_1_cry_0_Z));
    SLE \timeout_cnt[5]  (.D(timeout_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[5]));
    SLE \emflag_cnt[1]  (.D(emflag_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[1]));
    SLE \early_flags[123]  (.D(early_flags_7_fast_0[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[123]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[98]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[98]), .C(
        un10_early_flags[98]), .Y(late_flags_7_fast_0[98]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[27]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[27]), .C(
        un10_early_flags[27]), .Y(late_flags_7_fast_0[27]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[6]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[6]), .C(
        un10_early_flags[6]), .Y(late_flags_7_fast_0[6]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_18 (.A(
        early_flags_pmux_126_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[61]), .D(early_flags_Z[125]), .FCI(
        early_flags_pmux_126_1_1_co0_8), .S(
        early_flags_pmux_126_1_1_wmux_18_S_0), .Y(
        early_flags_pmux_126_1_1_y7_0), .FCO(
        early_flags_pmux_126_1_1_co1_8));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_23 (.A(
        un10_early_flags_2_0[16]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[20]), .Y(un10_early_flags[23]));
    SLE \late_flags[27]  (.D(late_flags_7_fast_0[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[27]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[2]), .D(
        late_flags_Z[66]), .FCI(VCC), .S(
        late_flags_pmux_63_1_0_wmux_S_0), .Y(
        late_flags_pmux_63_1_0_0_y0), .FCO(
        late_flags_pmux_63_1_0_0_co0));
    SLE \late_flags[60]  (.D(late_flags_7_fast_0[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[60]));
    CFG2 #( .INIT(4'hE) )  un1_bitalign_curr_state_13_1 (.A(
        early_flags_0_sqmuxa_1_Z), .B(bitalign_curr_state_Z[4]), .Y(
        un1_bitalign_curr_state_13_1_Z));
    CFG4 #( .INIT(16'h40C8) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNI7RVT2  (
        .A(bitalign_curr_state_Z[1]), .B(bitalign_curr_state149_1_Z), 
        .C(N_108), .D(N_63), .Y(i22_mux));
    CFG2 #( .INIT(4'h9) )  un1_bitalign_curr_state151 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state151_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_64 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_2_0[64]), .C(
        un10_early_flags_2_Z[8]), .Y(un10_early_flags[64]));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_0_wmux_8 (.A(
        early_flags_pmux_126_1_0_y0_3), .B(
        early_flags_pmux_126_1_0_0_y3), .C(
        early_flags_pmux_126_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_0_co0_3), .S(
        early_flags_pmux_126_1_0_wmux_8_S_0), .Y(
        early_flags_pmux_126_1_0_0_y9), .FCO(
        early_flags_pmux_126_1_0_co1_3));
    SLE \early_flags[2]  (.D(early_flags_7_fast_0[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[2]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_46 (.A(
        un10_early_flags_3_Z[46]), .B(tap_cnt_Z[6]), .C(
        un10_early_flags_1_Z[6]), .D(un10_early_flags_1_Z[40]), .Y(
        un10_early_flags[46]));
    SLE \late_flags[107]  (.D(late_flags_7_fast_0[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[107]));
    CFG2 #( .INIT(4'h8) )  
        \bitalign_curr_state_34_4_0_.un1_noearly_nolate_diff_start_valid  
        (.A(un2_noearly_nolate_diff_start_valid), .B(
        un1_early_late_diff_cry_7_Z), .Y(
        un1_noearly_nolate_diff_start_valid));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[122]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[122]), .C(
        un10_early_flags[122]), .Y(late_flags_7_fast_0[122]));
    SLE \early_flags[46]  (.D(early_flags_7_fast_0[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[46]));
    SLE \early_flags[47]  (.D(early_flags_7_fast_0[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[47]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[72]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[72]), .C(
        un10_early_flags[72]), .Y(late_flags_7_fast_0[72]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[118]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[118]), .C(
        un10_early_flags[118]), .Y(late_flags_7_fast_0[118]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_9 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_63_1_1_co1_3), .S(
        late_flags_pmux_63_1_1_wmux_9_S_0), .Y(
        late_flags_pmux_63_1_1_wmux_9_Y_0), .FCO(
        late_flags_pmux_63_1_1_co0_4));
    SLE \late_flags[77]  (.D(late_flags_7_fast_0[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[77]));
    SLE \early_late_diff[5]  (.D(early_late_diff_8[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[74]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[74]), .C(
        un10_early_flags[74]), .Y(early_flags_7_fast_0[74]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_7 (.A(
        late_flags_pmux_126_1_1_y7), .B(late_flags_pmux_126_1_1_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co1_2), .S(
        late_flags_pmux_126_1_1_wmux_7_S_0), .Y(
        late_flags_pmux_126_1_1_y0_3), .FCO(
        late_flags_pmux_126_1_1_co0_3));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_165  (.A(
        late_flags_Z[27]), .B(late_flags_Z[26]), .C(late_flags_Z[25]), 
        .D(late_flags_Z[24]), .Y(calc_done25_165));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[47]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[47]), .C(
        un10_early_flags[47]), .Y(late_flags_7_fast_0[47]));
    SLE \early_flags[41]  (.D(early_flags_7_fast_0[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[41]));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_114 (.A(tap_cnt_Z[3]), 
        .B(N_1499), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[114]));
    CFG4 #( .INIT(16'h8000) )  rx_BIT_ALGN_ERR (.A(timeout_cnt_Z[4]), 
        .B(timeout_cnt_Z[5]), .C(rx_BIT_ALGN_ERR_4_Z), .D(
        rx_BIT_ALGN_ERR_3_Z), .Y(BIT_ALGN_ERR_c));
    CFG2 #( .INIT(4'hE) )  un1_restart_trng_fg_10_0 (.A(
        un1_restart_trng_fg_10_sn_1), .B(tap_cnt_0_sqmuxa_1_Z), .Y(
        un1_restart_trng_fg_10_0_Z));
    CFG4 #( .INIT(16'hBFFF) )  \late_flags_7_i_o4[50]  (.A(
        tap_cnt_Z[0]), .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[48]), 
        .D(un10_early_flags_1_Z[48]), .Y(N_209));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_72 (.A(
        un10_early_flags_2_0[72]), .B(un10_early_flags_1_Z[0]), .C(
        un10_early_flags_1_Z[72]), .Y(un10_early_flags[72]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_16 (.A(
        early_flags_pmux_63_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[44]), .D(early_flags_Z[108]), .FCI(
        early_flags_pmux_63_1_1_co0_7), .S(
        early_flags_pmux_63_1_1_wmux_16_S_0), .Y(
        early_flags_pmux_63_1_1_y5_0), .FCO(
        early_flags_pmux_63_1_1_co1_7));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_14 (.A(
        early_flags_pmux_63_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[52]), .D(early_flags_Z[116]), .FCI(
        early_flags_pmux_63_1_1_co0_6), .S(
        early_flags_pmux_63_1_1_wmux_14_S_0), .Y(
        early_flags_pmux_63_1_1_y3_0), .FCO(
        early_flags_pmux_63_1_1_co1_6));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[3]), 
        .D(early_flags_Z[67]), .FCI(VCC), .S(
        early_flags_pmux_126_1_0_wmux_S_0), .Y(
        early_flags_pmux_126_1_0_0_y0), .FCO(
        early_flags_pmux_126_1_0_0_co0));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_168  (.A(
        late_flags_Z[47]), .B(late_flags_Z[46]), .C(late_flags_Z[45]), 
        .D(late_flags_Z[44]), .Y(calc_done25_168));
    SLE \late_flags[86]  (.D(late_flags_7_fast_0[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[86]));
    SLE \noearly_nolate_diff_nxt[5]  (.D(noearly_nolate_diff_nxt_8[5]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_5));
    SLE \early_late_diff[2]  (.D(early_late_diff_8[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[2]));
    SLE \late_flags[37]  (.D(late_flags_7_fast_0[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[37]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[23]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[23]), .C(
        un10_early_flags[23]), .Y(early_flags_7_fast_0[23]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_6 (.A(
        late_flags_pmux_63_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[56]), .D(late_flags_Z[120]), .FCI(
        late_flags_pmux_63_1_1_co0_2), .S(
        late_flags_pmux_63_1_1_wmux_6_S_0), .Y(
        late_flags_pmux_63_1_1_y7), .FCO(late_flags_pmux_63_1_1_co1_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[83]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[83]), .C(
        un10_early_flags[83]), .Y(early_flags_7_fast_0[83]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_4 (.A(
        un10_tapcnt_final_4), .B(early_late_diff_Z[4]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_3_Z), .S(
        un1_early_late_diff_cry_4_S_0), .Y(
        un1_early_late_diff_cry_4_Y_0), .FCO(
        un1_early_late_diff_cry_4_Z));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_4_0 (.A(
        emflag_cnt_Z[4]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[4]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_3), .S(
        noearly_nolate_diff_nxt_8[4]), .Y(
        noearly_nolate_diff_nxt_8_cry_4_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_4));
    CFG3 #( .INIT(8'h80) )  rx_BIT_ALGN_LOAD_0_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(tap_cnt_0_sqmuxa_2_0), .C(
        un1_bitalign_curr_state152_Z), .Y(rx_BIT_ALGN_LOAD_0_sqmuxa_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_184  (.A(
        late_flags_Z[119]), .B(late_flags_Z[118]), .C(
        late_flags_Z[117]), .D(late_flags_Z[116]), .Y(calc_done25_184));
    SLE rx_BIT_ALGN_MOVE (.D(rx_BIT_ALGN_MOVE_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE));
    SLE \late_flags[16]  (.D(late_flags_7_fast_0[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[16]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[12]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[12]), .C(
        un10_early_flags[12]), .Y(early_flags_7_fast_0[12]));
    CFG4 #( .INIT(16'hAAEA) )  un1_restart_trng_fg (.A(
        restart_trng_fg_i), .B(bitalign_curr_state148_2_Z), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        un1_restart_trng_fg_0));
    CFG4 #( .INIT(16'h8880) )  un1_early_late_diff_valid (.A(
        late_last_set_Z), .B(early_last_set_Z), .C(
        un2_early_late_diff_validlto7_2_Z), .D(
        un2_early_late_diff_validlt7), .Y(un1_early_late_diff_valid_Z));
    CFG4 #( .INIT(16'hFF13) )  un1_restart_trng_fg_6 (.A(
        bitalign_curr_state155), .B(tapcnt_final_upd_2_sqmuxa), .C(
        mv_dn_fg_Z), .D(restart_trng_fg_i), .Y(un1_restart_trng_fg_6_Z)
        );
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[104]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[104]), .C(
        un10_early_flags[104]), .Y(late_flags_7_fast_0[104]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[5]), 
        .D(early_flags_Z[69]), .FCI(early_flags_pmux_126_1_1_co1_4), 
        .S(early_flags_pmux_126_1_1_wmux_11_S_0), .Y(
        early_flags_pmux_126_1_1_y0_4), .FCO(
        early_flags_pmux_126_1_1_co0_5));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[63]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[63]), .C(
        un10_early_flags[63]), .Y(early_flags_7_fast_0[63]));
    SLE \early_flags[30]  (.D(early_flags_7_fast_0[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[30]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_135  (.A(
        early_flags_Z[107]), .B(early_flags_Z[106]), .C(
        early_flags_Z[105]), .D(early_flags_Z[104]), .Y(
        calc_done25_135));
    CFG2 #( .INIT(4'h8) )  mv_dn_fg_0_sqmuxa_i_a2_0 (.A(
        bitalign_curr_state148_Z), .B(un1_rx_BIT_ALGN_START), .Y(N_98));
    SLE \late_flags[55]  (.D(late_flags_7_fast_0[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[55]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[6]  (.A(VCC), .B(
        rst_cnt_Z[6]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[5]), .S(
        rst_cnt_s[6]), .Y(rst_cnt_cry_Y_1[6]), .FCO(rst_cnt_cry_Z[6]));
    CFG2 #( .INIT(4'h4) )  reset_dly_fg4_4 (.A(reset_dly_fg_Z), .B(
        rst_cnt_Z[9]), .Y(reset_dly_fg4_4_Z));
    SLE \early_flags[55]  (.D(early_flags_7_fast_0[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[55]));
    CFG4 #( .INIT(16'h353F) )  \bitalign_curr_state_34_4_0_.m50_1_1  (
        .A(bitalign_curr_state41_Z), .B(N_50), .C(
        bitalign_curr_state_Z[2]), .D(bitalign_curr_state_Z[0]), .Y(
        m50_1_1));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_4 (.A(
        early_flags_pmux_63_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[42]), .D(early_flags_Z[106]), .FCI(
        early_flags_pmux_63_1_0_co0_1), .S(
        early_flags_pmux_63_1_0_wmux_4_S_0), .Y(
        early_flags_pmux_63_1_0_0_y5), .FCO(
        early_flags_pmux_63_1_0_co1_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[98]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[98]), .C(
        un10_early_flags[98]), .Y(early_flags_7_fast_0[98]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[54]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[54]), .C(
        un10_early_flags[54]), .Y(late_flags_7_fast_0[54]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_104 (.A(
        un10_early_flags_1_Z[40]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[64]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[104]));
    SLE \tapcnt_final_upd[4]  (.D(tapcnt_final_upd_8[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[4]));
    SLE \late_flags[46]  (.D(late_flags_7_fast_0[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[46]));
    CFG4 #( .INIT(16'h10BA) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNI77PE2  (
        .A(bitalign_curr_state_Z[1]), .B(early_flags_dec[127]), .C(
        bitalign_curr_state89), .D(N_63), .Y(m82_1_1));
    ARI1 #( .INIT(20'h45500) )  early_late_diff_8_cry_0_0_cy (.A(VCC), 
        .B(un1_restart_trng_fg_5_0), .C(GND), .D(GND), .FCI(VCC), .S(
        early_late_diff_8_cry_0_0_cy_S_0), .Y(
        early_late_diff_8_cry_0_0_cy_Y_0), .FCO(
        early_late_diff_8_cry_0_0_cy_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_138  (.A(
        early_flags_Z[95]), .B(early_flags_Z[94]), .C(
        early_flags_Z[93]), .D(early_flags_Z[92]), .Y(calc_done25_138));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[95]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[95]), .C(
        un10_early_flags[95]), .Y(early_flags_7_fast_0[95]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_1_wmux_20 (.A(
        late_flags_pmux_126_1_1_y0_8), .B(late_flags_pmux_126_1_1_y3_0)
        , .C(late_flags_pmux_126_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co0_9), .S(
        late_flags_pmux_126_1_1_wmux_20_S_0), .Y(
        late_flags_pmux_126_1_1_y21), .FCO(
        late_flags_pmux_126_1_1_co1_9));
    CFG2 #( .INIT(4'h1) )  early_late_diff_0_sqmuxa_1_0 (.A(
        un1_tap_cnt_0_sqmuxa_6_0), .B(restart_trng_fg_i), .Y(
        early_late_diff_0_sqmuxa_1_0_Z));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_0 (.A(
        early_flags_pmux_126_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[35]), .D(early_flags_Z[99]), .FCI(
        early_flags_pmux_126_1_0_0_co0), .S(
        early_flags_pmux_126_1_0_wmux_0_S_0), .Y(
        early_flags_pmux_126_1_0_0_y1), .FCO(
        early_flags_pmux_126_1_0_0_co1));
    SLE \restart_edge_reg[3]  (.D(restart_edge_reg_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[3]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_14 (.A(
        late_flags_pmux_126_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[55]), .D(late_flags_Z[119]), .FCI(
        late_flags_pmux_126_1_0_co0_6), .S(
        late_flags_pmux_126_1_0_wmux_14_S_0), .Y(
        late_flags_pmux_126_1_0_y3_0), .FCO(
        late_flags_pmux_126_1_0_co1_6));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.calc_done26  (
        .A(calc_done25), .B(un1_tapcnt_final), .Y(calc_done26));
    CFG2 #( .INIT(4'hE) )  un1_early_flags_pmux_1 (.A(early_flags_pmux)
        , .B(late_flags_pmux), .Y(un1_early_flags_pmux_1_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_18 (.A(
        late_flags_pmux_126_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[61]), .D(late_flags_Z[125]), .FCI(
        late_flags_pmux_126_1_1_co0_8), .S(
        late_flags_pmux_126_1_1_wmux_18_S_0), .Y(
        late_flags_pmux_126_1_1_y7_0), .FCO(
        late_flags_pmux_126_1_1_co1_8));
    SLE \emflag_cnt[0]  (.D(emflag_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_18 (.A(
        late_flags_pmux_63_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[60]), .D(late_flags_Z[124]), .FCI(
        late_flags_pmux_63_1_1_co0_8), .S(
        late_flags_pmux_63_1_1_wmux_18_S_0), .Y(
        late_flags_pmux_63_1_1_y7_0), .FCO(
        late_flags_pmux_63_1_1_co1_8));
    SLE \noearly_nolate_diff_start[3]  (.D(
        noearly_nolate_diff_start_7[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_3));
    SLE \late_flags[81]  (.D(late_flags_7_fast_0[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[81]));
    CFG3 #( .INIT(8'hCE) )  \emflag_cnt_cry_cy_RNO[0]  (.A(
        bitalign_curr_state153_1_Z), .B(restart_trng_fg_i), .C(
        bitalign_curr_state_Z[1]), .Y(un1_restart_trng_fg_9_0_443_0));
    CFG4 #( .INIT(16'hAABA) )  rx_trng_done1_0_sqmuxa_i (.A(
        restart_trng_fg_i), .B(un1_bitalign_curr_state_16_1_Z), .C(
        N_52), .D(early_flags_0_sqmuxa_1_Z), .Y(
        rx_trng_done1_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI09J81[1]  (.A(early_val_Z[1])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[1]), .Y(
        early_val_RNI09J81_Z[1]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_237  (.A(
        calc_done25_183), .B(calc_done25_182), .C(calc_done25_181), .D(
        calc_done25_180), .Y(calc_done25_237));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[30]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[30]), .C(
        un10_early_flags[30]), .Y(late_flags_7_fast_0[30]));
    SLE \early_flags[60]  (.D(early_flags_7_fast_0[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[60]));
    ARI1 #( .INIT(20'h0F588) )  
        \bitalign_curr_state_34_4_0_.m74_2_1_1_wmux_0  (.A(
        m74_2_1_1_1_y0), .B(bitalign_curr_state_Z[1]), .C(N_29_i), .D(
        N_116_mux), .FCI(m74_2_1_1_1_co0), .S(m74_2_1_1_wmux_0_S_0), 
        .Y(N_75_0), .FCO(m74_2_1_1_1_co1));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_57 (.A(
        un10_early_flags_1_Z[9]), .B(tap_cnt_Z[6]), .C(
        un10_early_flags_1_Z[48]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[57]));
    CFG2 #( .INIT(4'h8) )  
        \bitalign_curr_state_34_4_0_.calc_done25_213  (.A(
        calc_done25_170), .B(calc_done25_171), .Y(calc_done25_213));
    CFG3 #( .INIT(8'h08) )  \bitalign_curr_state_34_4_0_.m110  (.A(
        bitalign_curr_state161_2_Z), .B(N_76_0), .C(
        bitalign_curr_state_Z[3]), .Y(N_130_mux));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_6 (.A(
        early_flags_pmux_126_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[59]), .D(early_flags_Z[123]), .FCI(
        early_flags_pmux_126_1_0_co0_2), .S(
        early_flags_pmux_126_1_0_wmux_6_S_0), .Y(
        early_flags_pmux_126_1_0_0_y7), .FCO(
        early_flags_pmux_126_1_0_co1_2));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[0]  (.A(
        no_early_no_late_val_end1_Z[0]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[0]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[0]));
    SLE \no_early_no_late_val_end2[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[0]));
    SLE \late_flags[65]  (.D(late_flags_7_fast_0[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[65]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[20]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[20]), .C(
        un10_early_flags[20]), .Y(late_flags_7_fast_0[20]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[116]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[116]), .C(
        un10_early_flags[116]), .Y(late_flags_7_fast_0[116]));
    CFG3 #( .INIT(8'hFB) )  early_cur_set_0_sqmuxa_i (.A(
        un1_tap_cnt_0_sqmuxa_6_0), .B(early_cur_set_0_sqmuxa_1_Z), .C(
        early_val_0_sqmuxa_1_0_Z), .Y(early_cur_set_0_sqmuxa_i_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_112 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_1_Z[48]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[112]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[29]), 
        .D(late_flags_Z[93]), .FCI(late_flags_pmux_126_1_1_co1_7), .S(
        late_flags_pmux_126_1_1_wmux_17_S_0), .Y(
        late_flags_pmux_126_1_1_y0_7), .FCO(
        late_flags_pmux_126_1_1_co0_8));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[25]), 
        .D(early_flags_Z[89]), .FCI(early_flags_pmux_126_1_1_co1_1), 
        .S(early_flags_pmux_126_1_1_wmux_5_S_0), .Y(
        early_flags_pmux_126_1_1_y0_2), .FCO(
        early_flags_pmux_126_1_1_co0_2));
    CFG2 #( .INIT(4'h8) )  rx_BIT_ALGN_ERR_3 (.A(timeout_cnt_Z[6]), .B(
        timeout_cnt_Z[7]), .Y(rx_BIT_ALGN_ERR_3_Z));
    SLE \late_flags[11]  (.D(late_flags_7_fast_0[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[11]));
    SLE \early_flags[32]  (.D(early_flags_7_fast_0[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[32]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIPPPT[3]  (.A(
        no_early_no_late_val_st1_Z[3]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[3]), .Y(
        un1_no_early_no_late_val_st1_1_1[3]));
    SLE \early_flags[7]  (.D(early_flags_7_fast_0[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[7]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_19 (.A(
        late_flags_pmux_63_1_0_y7_0), .B(late_flags_pmux_63_1_0_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co1_8), .S(
        late_flags_pmux_63_1_0_wmux_19_S_0), .Y(
        late_flags_pmux_63_1_0_y0_8), .FCO(
        late_flags_pmux_63_1_0_co0_9));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[11]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[11]), .C(
        un10_early_flags[11]), .Y(late_flags_7_fast_0[11]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_67 (.A(
        un10_early_flags_2_0[64]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_2_Z[67]), .Y(un10_early_flags[67]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[1]), 
        .D(early_flags_Z[65]), .FCI(VCC), .S(
        early_flags_pmux_126_1_1_wmux_S_0), .Y(
        early_flags_pmux_126_1_1_y0), .FCO(
        early_flags_pmux_126_1_1_co0));
    SLE \rst_cnt[7]  (.D(rst_cnt_s[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[7]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[103]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[103]), .C(
        un10_early_flags[103]), .Y(late_flags_7_fast_0[103]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[6]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[6]), .C(
        un10_early_flags[6]), .Y(early_flags_7_fast_0[6]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[12]), 
        .D(early_flags_Z[76]), .FCI(early_flags_pmux_63_1_1_co1_6), .S(
        early_flags_pmux_63_1_1_wmux_15_S_0), .Y(
        early_flags_pmux_63_1_1_y0_6), .FCO(
        early_flags_pmux_63_1_1_co0_7));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIHEIR[0]  (.A(
        late_val_Z[0]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[0]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIHEIR_0[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[74]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[74]), .C(
        un10_early_flags[74]), .Y(late_flags_7_fast_0[74]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[24]), 
        .D(late_flags_Z[88]), .FCI(late_flags_pmux_63_1_1_co1_1), .S(
        late_flags_pmux_63_1_1_wmux_5_S_0), .Y(
        late_flags_pmux_63_1_1_y0_2), .FCO(
        late_flags_pmux_63_1_1_co0_2));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_75 (.A(
        un10_early_flags_2_0[72]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[72]), .Y(un10_early_flags[75]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_121 (.A(
        un10_early_flags_1_Z[9]), .B(tap_cnt_Z[2]), .C(
        un10_early_flags_1_Z[48]), .D(un10_early_flags_2_Z[69]), .Y(
        un10_early_flags[121]));
    SLE \late_flags[41]  (.D(late_flags_7_fast_0[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[41]));
    SLE \early_flags[125]  (.D(early_flags_7_fast_0[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[125]));
    SLE \early_flags[48]  (.D(early_flags_7_fast_0[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[48]));
    SLE \late_flags[23]  (.D(late_flags_7_fast_0[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[23]));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_3_sqmuxa (.A(
        early_flags_1_sqmuxa_1_Z), .B(un1_rx_BIT_ALGN_START), .Y(
        tapcnt_final_upd_3_sqmuxa_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_99 (.A(
        un10_early_flags_1_Z[3]), .B(un10_early_flags_2_0[96]), .C(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[99]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_4_0 (.A(
        emflag_cnt_Z[4]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[4]), .D(GND), .FCI(early_late_diff_8_cry_3), .S(
        early_late_diff_8[4]), .Y(early_late_diff_8_cry_4_0_Y_0), .FCO(
        early_late_diff_8_cry_4));
    SLE \late_flags[96]  (.D(late_flags_7_fast_0[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[96]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[40]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[40]), .C(
        un10_early_flags[40]), .Y(late_flags_7_fast_0[40]));
    CFG4 #( .INIT(16'h0040) )  bitalign_curr_state_0_sqmuxa_10_0_a2 (
        .A(un1_retrain_adj_tap_i), .B(un1_rx_BIT_ALGN_START), .C(
        bitalign_curr_state148_Z), .D(bitalign_curr_state12_Z), .Y(
        bitalign_curr_state_0_sqmuxa_10));
    SLE \early_flags[70]  (.D(early_flags_7_fast_0[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[70]));
    SLE \early_flags[62]  (.D(early_flags_7_fast_0[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[62]));
    SLE \early_flags[117]  (.D(early_flags_7_fast_0[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[117]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_56 (.A(
        un10_early_flags_1_Z[32]), .B(tap_cnt_Z[6]), .C(
        un10_early_flags_1_Z[24]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[56]));
    SLE early_last_set (.D(early_last_set_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_last_set_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(early_last_set_Z)
        );
    CFG3 #( .INIT(8'hAB) )  tapcnt_final_upd_0_sqmuxa_i (.A(
        restart_trng_fg_i), .B(un1_bitalign_curr_state_13_1_Z), .C(
        un1_bitalign_curr_state_14_1_0_Z), .Y(
        tapcnt_final_upd_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[124]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[124]), .C(
        un10_early_flags[124]), .Y(late_flags_7_fast_0[124]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_150  (.A(
        early_flags_Z[47]), .B(early_flags_Z[46]), .C(
        early_flags_Z[45]), .D(early_flags_Z[44]), .Y(calc_done25_150));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_0_0 (.A(
        emflag_cnt_Z[0]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[0]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Z), .S(
        noearly_nolate_diff_nxt_8[0]), .Y(
        noearly_nolate_diff_nxt_8_cry_0_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_0));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_0_wmux_20 (.A(
        early_flags_pmux_126_1_0_y0_8), .B(
        early_flags_pmux_126_1_0_y3_0), .C(
        early_flags_pmux_126_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_0_co0_9), .S(
        early_flags_pmux_126_1_0_wmux_20_S_0), .Y(
        early_flags_pmux_126_1_0_0_y21), .FCO(
        early_flags_pmux_126_1_0_co1_9));
    CFG2 #( .INIT(4'h7) )  un10_early_flags_17_1_i (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[0]), .Y(N_1498));
    CFG4 #( .INIT(16'hA5EC) )  \tapcnt_final_13_1[0]  (.A(
        tapcnt_final_13_1_1_0_Z[0]), .B(tapcnt_final_13_Z[1]), .C(
        tapcnt_final_13_m0s2_0), .D(un1_tapcnt_final_0_sqmuxa_Z), .Y(
        tapcnt_final_13_1_Z[0]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_102 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[96]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_2_Z[6]), .Y(
        un10_early_flags[102]));
    SLE rx_err (.D(N_1392), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_err_0_sqmuxa_1_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_err_Z));
    SLE \early_flags[85]  (.D(early_flags_7_fast_0[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[85]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[65]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[65]), .C(
        un10_early_flags[65]), .Y(late_flags_7_fast_0[65]));
    CFG1 #( .INIT(2'h1) )  \cnt_RNO[0]  (.A(CO0_0), .Y(CO0_0_i));
    SLE bit_align_start (.D(N_1439_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        bit_align_done_0_sqmuxa_3_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        bit_align_start_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_5 (.A(
        un10_tapcnt_final_5), .B(early_late_diff_Z[5]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_4_Z), .S(
        un1_early_late_diff_cry_5_S_0), .Y(
        un1_early_late_diff_cry_5_Y_0), .FCO(
        un1_early_late_diff_cry_5_Z));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_66 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[6]), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[66]));
    SLE \late_flags[73]  (.D(late_flags_7_fast_0[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[73]));
    SLE \early_flags[23]  (.D(early_flags_7_fast_0[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[23]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[4]  (.A(
        tapcnt_final_Z[4]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[4]), .Y(
        tapcnt_final_13_Z[4]));
    SLE \rst_cnt[0]  (.D(rst_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[0]));
    SLE \late_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[3])
        );
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_6 (.A(
        late_flags_pmux_126_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[57]), .D(late_flags_Z[121]), .FCI(
        late_flags_pmux_126_1_1_co0_2), .S(
        late_flags_pmux_126_1_1_wmux_6_S_0), .Y(
        late_flags_pmux_126_1_1_y7), .FCO(
        late_flags_pmux_126_1_1_co1_2));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_176  (.A(
        late_flags_Z[87]), .B(late_flags_Z[86]), .C(late_flags_Z[85]), 
        .D(late_flags_Z[84]), .Y(calc_done25_176));
    CFG2 #( .INIT(4'h2) )  
        \bitalign_curr_state_34_4_0_.un1_tapcnt_final  (.A(un34), .B(
        un16_tapcnt_final_cry_7_Z), .Y(un1_tapcnt_final));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_7 (.A(
        un16_tapcnt_final_7), .B(early_late_diff_Z[7]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_6_Z), .S(
        un1_early_late_diff_1_cry_7_S_0), .Y(
        un1_early_late_diff_1_cry_7_Y_0), .FCO(
        un1_early_late_diff_1_cry_7_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[17]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[17]), .C(
        un10_early_flags[17]), .Y(early_flags_7_fast_0[17]));
    ARI1 #( .INIT(20'h472D8) )  \tap_cnt_RNO_0[6]  (.A(
        un1_tap_cnt_0_sqmuxa_14_0_0[1]), .B(N_60), .C(tap_cnt_Z[6]), 
        .D(tapcnt_final_Z[6]), .FCI(tap_cnt_17_i_m2_cry_5), .S(N_74), 
        .Y(tap_cnt_RNO_0_Y_0[6]), .FCO(tap_cnt_RNO_0_FCO_0[6]));
    CFG3 #( .INIT(8'h04) )  early_last_set_2_sqmuxa (.A(
        restart_trng_fg_i), .B(early_val_0_sqmuxa_1_0_Z), .C(
        early_flags_pmux), .Y(early_last_set_2_sqmuxa_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_10 (.A(
        early_flags_pmux_63_1_0_0_y21), .B(
        early_flags_pmux_63_1_0_0_y9), .C(emflag_cnt_Z[2]), .D(VCC), 
        .FCI(early_flags_pmux_63_1_0_co0_4), .S(
        early_flags_pmux_63_1_0_wmux_10_S_0), .Y(
        early_flags_pmux_63_1_0_wmux_10_Y_0), .FCO(
        early_flags_pmux_63_1_0_co1_4));
    CFG4 #( .INIT(16'h0007) )  rx_BIT_ALGN_MOVE_0_sqmuxa_2_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(
        rx_BIT_ALGN_MOVE_0_sqmuxa_0_Z), .C(
        un1_early_flags_1_sqmuxa_1_Z), .D(
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), .Y(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_1_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[119]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[119]), .C(
        un10_early_flags[119]), .Y(early_flags_7_fast_0[119]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[4]  (.A(VCC), .B(
        rst_cnt_Z[4]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[3]), .S(
        rst_cnt_s[4]), .Y(rst_cnt_cry_Y_1[4]), .FCO(rst_cnt_cry_Z[4]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_19 (.A(
        early_flags_pmux_126_1_1_y7_0), .B(
        early_flags_pmux_126_1_1_y5_0), .C(emflag_cnt_Z[4]), .D(
        emflag_cnt_Z[3]), .FCI(early_flags_pmux_126_1_1_co1_8), .S(
        early_flags_pmux_126_1_1_wmux_19_S_0), .Y(
        early_flags_pmux_126_1_1_y0_8), .FCO(
        early_flags_pmux_126_1_1_co0_9));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_2 (.A(
        early_flags_pmux_126_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[51]), .D(early_flags_Z[115]), .FCI(
        early_flags_pmux_126_1_0_co0_0), .S(
        early_flags_pmux_126_1_0_wmux_2_S_0), .Y(
        early_flags_pmux_126_1_0_0_y3), .FCO(
        early_flags_pmux_126_1_0_co1_0));
    SLE \late_flags[33]  (.D(late_flags_7_fast_0[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[33]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[93]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[93]), .C(
        un10_early_flags[93]), .Y(early_flags_7_fast_0[93]));
    SLE \early_flags[72]  (.D(early_flags_7_fast_0[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[72]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_187  (.A(
        late_flags_Z[123]), .B(late_flags_Z[122]), .C(
        late_flags_Z[121]), .D(late_flags_Z[120]), .Y(calc_done25_187));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[38]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[38]), .C(
        un10_early_flags[38]), .Y(late_flags_7_fast_0[38]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_78 (.A(
        un10_early_flags_1_Z[72]), .B(un10_early_flags_1_Z[6]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_3_Z[46]), .Y(
        un10_early_flags[78]));
    SLE \bitalign_curr_state[1]  (.D(bitalign_curr_state_34[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[13]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[13]), .C(
        un10_early_flags[13]), .Y(late_flags_7_fast_0[13]));
    SLE \late_flags[91]  (.D(late_flags_7_fast_0[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[91]));
    SLE \restart_edge_reg[0]  (.D(Restart_trng_edge_det_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[0]));
    SLE \early_flags[95]  (.D(early_flags_7_fast_0[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[95]));
    CFG2 #( .INIT(4'h8) )  emflag_cnt_0_sqmuxa_1 (.A(
        bitalign_curr_state163_Z), .B(bit_align_dly_done_Z), .Y(
        emflag_cnt_0_sqmuxa_1_Z));
    CFG4 #( .INIT(16'h5150) )  rx_BIT_ALGN_LOAD_9_iv (.A(
        restart_trng_fg_i), .B(rx_err_Z), .C(un1_tap_cnt_0_sqmuxa_6_0), 
        .D(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .Y(rx_BIT_ALGN_LOAD_9)
        );
    SLE \rst_cnt[4]  (.D(rst_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[78]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[78]), .C(
        un10_early_flags[78]), .Y(early_flags_7_fast_0[78]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[28]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[28]), .C(
        un10_early_flags[28]), .Y(late_flags_7_fast_0[28]));
    CFG2 #( .INIT(4'h2) )  bitalign_curr_state154 (.A(
        bitalign_curr_state154_3_Z), .B(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state154_Z));
    CFG4 #( .INIT(16'h00CD) )  \bitalign_curr_state_34_4_0_.m67  (.A(
        m67_1), .B(m66_1), .C(bitalign_curr_state_Z[3]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[1]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[123]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[123]), .C(
        un10_early_flags[123]), .Y(late_flags_7_fast_0[123]));
    SLE \emflag_cnt[6]  (.D(emflag_cnt_s_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[6]));
    SLE \late_flags[120]  (.D(late_flags_7_fast_0[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[120]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_76_2_0 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[5]), .Y(
        un10_early_flags_2_0[76]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[75]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[75]), .C(
        un10_early_flags[75]), .Y(early_flags_7_fast_0[75]));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_2 (.A(
        tapcnt_final_upd_Z[2]), .B(tapcnt_final_Z[2]), .C(tap_cnt_Z[2])
        , .D(N_1416), .Y(bitalign_curr_state61_2_Z));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[6]  (.A(N_74), .B(N_63_0), .Y(
        N_1496_i));
    SLE \late_flags[8]  (.D(late_flags_7_fast_0[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[8]));
    SLE \rst_cnt[2]  (.D(rst_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[2]));
    CFG3 #( .INIT(8'h20) )  rx_err_1_sqmuxa (.A(
        bitalign_curr_state162_Z), .B(un1_calc_done25_7_i), .C(
        early_flags_dec[127]), .Y(rx_err_1_sqmuxa_Z));
    SLE \no_early_no_late_val_end2[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[6]));
    SLE \early_flags[0]  (.D(early_flags_7_fast_0[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[0]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_226  (.A(
        calc_done25_139), .B(calc_done25_138), .C(calc_done25_137), .D(
        calc_done25_136), .Y(calc_done25_226));
    SLE calc_done (.D(N_1431_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(calc_done_0_sqmuxa_2_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(calc_done_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_83 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[0]), .Y(
        un10_early_flags[83]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_140  (.A(
        early_flags_Z[71]), .B(early_flags_Z[70]), .C(
        early_flags_Z[69]), .D(early_flags_Z[68]), .Y(calc_done25_140));
    SLE \early_flags[110]  (.D(early_flags_7_fast_0[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[110]));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[5]  (.A(N_75), .B(N_63_0), .Y(
        N_1497_i));
    SLE \noearly_nolate_diff_nxt[2]  (.D(noearly_nolate_diff_nxt_8[2]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_2));
    CFG3 #( .INIT(8'hF4) )  un1_bitalign_curr_state148_8_0 (.A(
        bit_align_dly_done_Z), .B(bitalign_curr_state163_Z), .C(
        timeout_cnt_1_sqmuxa_Z), .Y(un1_bitalign_curr_state148_8_0_Z));
    SLE \no_early_no_late_val_end1[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[2]));
    SLE \no_early_no_late_val_end2[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[48]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[48]), .C(
        un10_early_flags[48]), .Y(late_flags_7_fast_0[48]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_12 (.A(
        early_flags_pmux_126_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[39]), .D(early_flags_Z[103]), .FCI(
        early_flags_pmux_126_1_0_co0_5), .S(
        early_flags_pmux_126_1_0_wmux_12_S_0), .Y(
        early_flags_pmux_126_1_0_y1_0), .FCO(
        early_flags_pmux_126_1_0_co1_5));
    SLE \late_flags[29]  (.D(late_flags_7_fast_0[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[29]));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.m34  (.A(
        early_flags_pmux), .B(early_cur_set_Z), .Y(N_35));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_123 (.A(
        un10_early_flags_1_Z[24]), .B(tap_cnt_Z[2]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[96]), .Y(
        un10_early_flags[123]));
    SLE \no_early_no_late_val_st1[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[81]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[81]), .C(
        un10_early_flags[81]), .Y(late_flags_7_fast_0[81]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[119]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[119]), .C(
        un10_early_flags[119]), .Y(late_flags_7_fast_0[119]));
    ARI1 #( .INIT(20'h4B4AA) )  \tapcnt_final_13_RNO[6]  (.A(
        un1_bitalign_curr_state169_12_sn), .B(early_val_Z[6]), .C(
        tapcnt_final_3_sqmuxa_Z), .D(tapcnt_final_13_m1_axb_6_1), .FCI(
        tapcnt_final_13_m1_cry_5), .S(tapcnt_final_13_m1[6]), .Y(
        tapcnt_final_13_RNO_Y_0[6]), .FCO(tapcnt_final_13_RNO_FCO_0[6])
        );
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_174  (.A(
        late_flags_Z[55]), .B(late_flags_Z[54]), .C(late_flags_Z[53]), 
        .D(late_flags_Z[52]), .Y(calc_done25_174));
    CFG2 #( .INIT(4'h8) )  early_val_0_sqmuxa_1_0 (.A(
        bitalign_curr_state160_Z), .B(early_cur_set_Z), .Y(
        early_val_0_sqmuxa_1_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[67]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[67]), .C(
        un10_early_flags[67]), .Y(late_flags_7_fast_0[67]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_248  (.A(
        calc_done25_227), .B(calc_done25_226), .C(calc_done25_225), .D(
        calc_done25_224), .Y(calc_done25_248));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_71 (.A(tap_cnt_Z[6]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[71]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[19]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[19]), .C(
        un10_early_flags[19]), .Y(early_flags_7_fast_0[19]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_6 (.A(late_val_Z[6])
        , .B(early_val_Z[6]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_5_Z), .S(tapcnt_final27_cry_6_S_0), .Y(
        tapcnt_final27_cry_6_Y_0), .FCO(tapcnt_final27));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_39 (.A(
        un10_early_flags_2_0[32]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[36]), .Y(un10_early_flags[39]));
    SLE \early_flags[4]  (.D(early_flags_7_fast_0[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[4]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_155  (.A(
        early_flags_Z[27]), .B(early_flags_Z[26]), .C(
        early_flags_Z[25]), .D(early_flags_Z[24]), .Y(calc_done25_155));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[36]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[36]), .C(
        un10_early_flags[36]), .Y(early_flags_7_fast_0[36]));
    SLE \late_flags[79]  (.D(late_flags_7_fast_0[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[79]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_2 (.A(
        un10_tapcnt_final_2), .B(early_late_diff_Z[2]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_1_Z), .S(
        un1_early_late_diff_cry_2_S_0), .Y(
        un1_early_late_diff_cry_2_Y_0), .FCO(
        un1_early_late_diff_cry_2_Z));
    CFG4 #( .INIT(16'h30A3) )  un1_bitalign_curr_state148_2 (.A(
        bitalign_curr_state152_1_Z), .B(un1_bitalign_curr_state_14_1_Z)
        , .C(bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[2]), 
        .Y(un1_bitalign_curr_state148_2_Z));
    SLE \no_early_no_late_val_end2[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[1]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_1 (.A(
        un10_tapcnt_final_1), .B(early_late_diff_Z[1]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_0_Z), .S(
        un1_early_late_diff_cry_1_S_0), .Y(
        un1_early_late_diff_cry_1_Y_0), .FCO(
        un1_early_late_diff_cry_1_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[2]), 
        .D(early_flags_Z[66]), .FCI(VCC), .S(
        early_flags_pmux_63_1_0_wmux_S_0), .Y(
        early_flags_pmux_63_1_0_0_y0), .FCO(
        early_flags_pmux_63_1_0_0_co0));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_158  (.A(
        early_flags_Z[7]), .B(early_flags_Z[6]), .C(early_flags_Z[5]), 
        .D(early_flags_Z[4]), .Y(calc_done25_158));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_0_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(un10_early_flags_2_0[0])
        );
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[40]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[40]), .C(
        un10_early_flags[40]), .Y(early_flags_7_fast_0[40]));
    CFG4 #( .INIT(16'hFFFE) )  un1_bitalign_curr_state_1_sqmuxa_6 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_Z), .B(
        early_flags_0_sqmuxa_Z), .C(bitalign_curr_state_1_sqmuxa_4_Z), 
        .D(bit_align_done_0_sqmuxa_2_Z), .Y(
        un1_bitalign_curr_state_1_sqmuxa_6_i_0));
    CFG4 #( .INIT(16'h4CCC) )  timeout_cnt_1_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state154_Z), 
        .C(rx_err_Z), .D(calc_done_Z), .Y(timeout_cnt_1_sqmuxa_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_29 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_2_0[28]), .C(
        un10_early_flags_1_Z[5]), .Y(un10_early_flags[29]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[7]  (.A(VCC), .B(
        rst_cnt_Z[7]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[6]), .S(
        rst_cnt_s[7]), .Y(rst_cnt_cry_Y_1[7]), .FCO(rst_cnt_cry_Z[7]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[0]), .D(
        late_flags_Z[64]), .FCI(VCC), .S(
        late_flags_pmux_63_1_1_wmux_S_0), .Y(late_flags_pmux_63_1_1_y0)
        , .FCO(late_flags_pmux_63_1_1_co0));
    CFG3 #( .INIT(8'h80) )  bitalign_curr_state_0_sqmuxa_9 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state155), .C(
        bitalign_curr_state61), .Y(bitalign_curr_state_0_sqmuxa_9_Z));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_1_wmux_8 (.A(
        early_flags_pmux_63_1_1_y0_3), .B(early_flags_pmux_63_1_1_y3), 
        .C(early_flags_pmux_63_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co0_3), .S(
        early_flags_pmux_63_1_1_wmux_8_S_0), .Y(
        early_flags_pmux_63_1_1_y9), .FCO(
        early_flags_pmux_63_1_1_co1_3));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_19 (.A(
        late_flags_pmux_63_1_1_y7_0), .B(late_flags_pmux_63_1_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co1_8), .S(
        late_flags_pmux_63_1_1_wmux_19_S_0), .Y(
        late_flags_pmux_63_1_1_y0_8), .FCO(
        late_flags_pmux_63_1_1_co0_9));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[19]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[19]), .C(
        un10_early_flags[19]), .Y(late_flags_7_fast_0[19]));
    SLE \late_flags[39]  (.D(late_flags_7_fast_0[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[39]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_7 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[7]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_70 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[64]), .C(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[70]));
    SLE \late_flags[88]  (.D(late_flags_7_fast_0[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[88]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_16_1 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[16]));
    SLE \late_flags[52]  (.D(late_flags_7_fast_0[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[52]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_224  (.A(
        calc_done25_131), .B(calc_done25_130), .C(calc_done25_129), .D(
        calc_done25_128), .Y(calc_done25_224));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_6 (.A(
        un16_tapcnt_final_6), .B(early_late_diff_Z[6]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_5_Z), .S(
        un1_early_late_diff_1_cry_6_S_0), .Y(
        un1_early_late_diff_1_cry_6_Y_0), .FCO(
        un1_early_late_diff_1_cry_6_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[54]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[54]), .C(
        un10_early_flags[54]), .Y(early_flags_7_fast_0[54]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_5_0 (.A(
        emflag_cnt_Z[5]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[5]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_4), .S(
        noearly_nolate_diff_nxt_8[5]), .Y(
        noearly_nolate_diff_nxt_8_cry_5_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_5));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_2 (.A(
        un10_tapcnt_final_2), .B(un16_tapcnt_final_2), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_1_Z), .S(
        un10_tapcnt_final_cry_2_S_0), .Y(un10_tapcnt_final_cry_2_Y_0), 
        .FCO(un10_tapcnt_final_cry_2_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_36_1 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[36]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_2_0 (.A(
        emflag_cnt_Z[2]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[2]), .D(GND), .FCI(early_late_diff_8_cry_1), .S(
        early_late_diff_8[2]), .Y(early_late_diff_8_cry_2_0_Y_0), .FCO(
        early_late_diff_8_cry_2));
    SLE \late_flags[104]  (.D(late_flags_7_fast_0[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[104]));
    SLE \early_flags[122]  (.D(early_flags_7_fast_0[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[122]));
    SLE bit_align_dly_done (.D(bit_align_dly_done_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        bit_align_dly_done_0_sqmuxa_1_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bit_align_dly_done_Z));
    SLE \late_flags[0]  (.D(late_flags_7_fast_0[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[0]));
    SLE \restart_reg[1]  (.D(restart_reg_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_reg_Z[1]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_6_0 (
        .A(emflag_cnt_Z[6]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[6]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_5), .S(
        noearly_nolate_diff_start_7[6]), .Y(
        noearly_nolate_diff_start_7_cry_6_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_6));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_13 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[3]), .C(un10_early_flags_1_Z[5]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[13]));
    SLE \late_flags[18]  (.D(late_flags_7_fast_0[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[18]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_4 (.A(
        late_flags_pmux_63_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[40]), .D(late_flags_Z[104]), .FCI(
        late_flags_pmux_63_1_1_co0_1), .S(
        late_flags_pmux_63_1_1_wmux_4_S_0), .Y(
        late_flags_pmux_63_1_1_y5), .FCO(late_flags_pmux_63_1_1_co1_1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[83]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[83]), .C(
        un10_early_flags[83]), .Y(late_flags_7_fast_0[83]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[116]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[116]), .C(
        un10_early_flags[116]), .Y(early_flags_7_fast_0[116]));
    CFG2 #( .INIT(4'h1) )  bitalign_curr_state148_2 (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[4]), .Y(
        bitalign_curr_state148_2_Z));
    CFG4 #( .INIT(16'hCCDF) )  rx_err_0_sqmuxa_1_i (.A(
        bitalign_curr_state162_Z), .B(restart_trng_fg_i), .C(
        un1_calc_done25_7_i), .D(un1_bitalign_curr_state148_9_2_Z), .Y(
        rx_err_0_sqmuxa_1_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[73]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[73]), .C(
        un10_early_flags[73]), .Y(early_flags_7_fast_0[73]));
    CFG4 #( .INIT(16'hFFFE) )  \bitalign_curr_state_34_4_0_.un34lto7  
        (.A(un16_tapcnt_final_4), .B(un16_tapcnt_final_5), .C(
        un34lto7_4), .D(un34lto7_3), .Y(un34));
    CFG2 #( .INIT(4'hE) )  \un1_tap_cnt_0_sqmuxa_14_0_o2_0[1]  (.A(
        un1_bitalign_curr_state_1_sqmuxa_2_i_0), .B(
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), .Y(N_82));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_1_0 (
        .A(emflag_cnt_Z[1]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[1]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_0), .S(
        noearly_nolate_diff_start_7[1]), .Y(
        noearly_nolate_diff_start_7_cry_1_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_1));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_6 (.A(
        early_flags_pmux_63_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[58]), .D(early_flags_Z[122]), .FCI(
        early_flags_pmux_63_1_0_co0_2), .S(
        early_flags_pmux_63_1_0_wmux_6_S_0), .Y(
        early_flags_pmux_63_1_0_0_y7), .FCO(
        early_flags_pmux_63_1_0_co1_2));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_9 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_63_1_0_co1_3), .S(
        late_flags_pmux_63_1_0_wmux_9_S_0), .Y(
        late_flags_pmux_63_1_0_wmux_9_Y_0), .FCO(
        late_flags_pmux_63_1_0_co0_4));
    SLE \early_flags[54]  (.D(early_flags_7_fast_0[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[54]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_4 (.A(
        un16_tapcnt_final_4), .B(un10_tapcnt_final_4), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_3_Z), .S(
        un16_tapcnt_final_cry_4_S_0), .Y(un16_tapcnt_final_cry_4_Y_0), 
        .FCO(un16_tapcnt_final_cry_4_Z));
    CFG4 #( .INIT(16'hFEFF) )  un1_bitalign_curr_state148_9_2 (.A(
        rx_trng_done_1_sqmuxa_Z), .B(timeout_cnt_1_sqmuxa_Z), .C(
        un1_bitalign_curr_state148_8_1_Z), .D(
        un1_bitalign_curr_state148_5_Z), .Y(
        un1_bitalign_curr_state148_9_2_Z));
    SLE \early_flags[43]  (.D(early_flags_7_fast_0[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[43]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_232  (.A(
        calc_done25_163), .B(calc_done25_162), .C(calc_done25_161), .D(
        calc_done25_160), .Y(calc_done25_232));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[44]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[44]), .C(
        un10_early_flags[44]), .Y(early_flags_7_fast_0[44]));
    SLE \late_flags[48]  (.D(late_flags_7_fast_0[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[48]));
    SLE \late_flags[62]  (.D(late_flags_7_fast_0[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[62]));
    CFG4 #( .INIT(16'h083B) )  \bitalign_curr_state_34_4_0_.m86_1  (.A(
        bitalign_curr_state161_2_Z), .B(bitalign_curr_state_Z[4]), .C(
        N_76_0), .D(N_75_0), .Y(m86_1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[16]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[16]), .C(
        un10_early_flags[16]), .Y(late_flags_7_fast_0[16]));
    SLE \late_flags[123]  (.D(late_flags_7_fast_0[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[123]));
    SLE \late_flags[109]  (.D(late_flags_7_fast_0[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[109]));
    SLE \early_late_diff[3]  (.D(early_late_diff_8[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[3]));
    CFG4 #( .INIT(16'h4C7F) )  \bitalign_curr_state_34_4_0_.m101_1_1  
        (.A(bitalign_curr_state161_2_Z), .B(bitalign_curr_state_Z[4]), 
        .C(N_94), .D(N_92), .Y(m101_1_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[109]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[109]), .C(
        un10_early_flags[109]), .Y(early_flags_7_fast_0[109]));
    SLE \early_late_diff[6]  (.D(early_late_diff_8[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[6]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_145  (.A(
        early_flags_Z[51]), .B(early_flags_Z[50]), .C(
        early_flags_Z[49]), .D(early_flags_Z[48]), .Y(calc_done25_145));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_1 (.A(
        tapcnt_final_upd_Z[1]), .B(tapcnt_final_Z[1]), .C(tap_cnt_Z[1])
        , .D(N_1416), .Y(bitalign_curr_state61_1_Z));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_16 (.A(
        early_flags_pmux_126_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[47]), .D(early_flags_Z[111]), .FCI(
        early_flags_pmux_126_1_0_co0_7), .S(
        early_flags_pmux_126_1_0_wmux_16_S_0), .Y(
        early_flags_pmux_126_1_0_y5_0), .FCO(
        early_flags_pmux_126_1_0_co1_7));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_111 (.A(
        un10_early_flags_1_Z[96]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[111]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[91]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[91]), .C(
        un10_early_flags[91]), .Y(late_flags_7_fast_0[91]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[115]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[115]), .C(
        un10_early_flags[115]), .Y(early_flags_7_fast_0[115]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_6 (.A(
        late_flags_pmux_63_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[58]), .D(late_flags_Z[122]), .FCI(
        late_flags_pmux_63_1_0_co0_2), .S(
        late_flags_pmux_63_1_0_wmux_6_S_0), .Y(
        late_flags_pmux_63_1_0_0_y7), .FCO(
        late_flags_pmux_63_1_0_co1_2));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[100]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[100]), .C(
        un10_early_flags[100]), .Y(late_flags_7_fast_0[100]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[114]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[114]), .C(
        un10_early_flags[114]), .Y(early_flags_7_fast_0[114]));
    CFG4 #( .INIT(16'h0013) )  bit_align_done_0_sqmuxa_3_1 (.A(
        bitalign_curr_state161_2_Z), .B(
        bitalign_curr_state_1_sqmuxa_4_Z), .C(
        bit_align_dly_done_0_sqmuxa_1_0_Z), .D(restart_trng_fg_i), .Y(
        bit_align_done_0_sqmuxa_3_1_Z));
    SLE \late_flags[121]  (.D(late_flags_7_fast_0[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[121]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[5]  (.A(VCC), .B(
        rst_cnt_Z[5]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[4]), .S(
        rst_cnt_s[5]), .Y(rst_cnt_cry_Y_1[5]), .FCO(rst_cnt_cry_Z[5]));
    SLE \tapcnt_final_upd[2]  (.D(tapcnt_final_upd_8_cry_2_0_Y_0), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[2]));
    SLE sig_rx_BIT_ALGN_CLR_FLGS (.D(sig_rx_BIT_ALGN_CLR_FLGS_11), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(sig_rx_BIT_ALGN_CLR_FLGS_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_63_1_0_co1_3), .S(
        early_flags_pmux_63_1_0_wmux_9_S_0), .Y(
        early_flags_pmux_63_1_0_wmux_9_Y_0), .FCO(
        early_flags_pmux_63_1_0_co0_4));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_10 (.A(
        early_flags_pmux_126_1_1_y21), .B(early_flags_pmux_126_1_1_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_126_1_1_co0_4), .S(
        early_flags_pmux_126_1_1_wmux_10_S_0), .Y(
        early_flags_pmux_126_1_1_wmux_10_Y_0), .FCO(
        early_flags_pmux_126_1_1_co1_4));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_148  (.A(
        early_flags_Z[39]), .B(early_flags_Z[38]), .C(
        early_flags_Z[37]), .D(early_flags_Z[36]), .Y(calc_done25_148));
    CFG3 #( .INIT(8'hFE) )  un1_tapcnt_final_0_sqmuxa (.A(
        tapcnt_final_5_sqmuxa), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .Y(un1_tapcnt_final_0_sqmuxa_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_s[9]  (.A(VCC), .B(
        rst_cnt_Z[9]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[8]), .S(
        rst_cnt_s_Z[9]), .Y(rst_cnt_s_Y_1[9]), .FCO(rst_cnt_s_FCO_1[9])
        );
    SLE \late_flags[84]  (.D(late_flags_7_fast_0[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[84]));
    CFG3 #( .INIT(8'h04) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state155  (.A(
        un1_bitalign_curr_state_15_1_Z), .B(bitalign_curr_state155_1), 
        .C(bitalign_curr_state_Z[3]), .Y(bitalign_curr_state155));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[117]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[117]), .C(
        un10_early_flags[117]), .Y(late_flags_7_fast_0[117]));
    SLE \late_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[4])
        );
    SLE \early_flags[56]  (.D(early_flags_7_fast_0[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[56]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_129  (.A(
        early_flags_Z[115]), .B(early_flags_Z[114]), .C(
        early_flags_Z[113]), .D(early_flags_Z[112]), .Y(
        calc_done25_129));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[60]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[60]), .C(
        un10_early_flags[60]), .Y(late_flags_7_fast_0[60]));
    SLE \early_flags[57]  (.D(early_flags_7_fast_0[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[57]));
    CFG3 #( .INIT(8'h02) )  bitalign_curr_state149 (.A(
        bitalign_curr_state149_1_Z), .B(un1_bitalign_curr_state_14_1_Z)
        , .C(bitalign_curr_state_Z[4]), .Y(bitalign_curr_state149_Z));
    CFG4 #( .INIT(16'h00A8) )  calc_done_RNO (.A(
        bitalign_curr_state_Z[4]), .B(early_flags_dec[127]), .C(
        un1_calc_done25_7_i), .D(restart_trng_fg_i), .Y(N_1431_i));
    CFG3 #( .INIT(8'h5D) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state159_RNIPFGK  (
        .A(early_late_diff_0_sqmuxa_1_0_Z), .B(bitalign_curr_state159), 
        .C(un1_early_flags_pmux_1_Z), .Y(
        no_early_no_late_val_end1_0_sqmuxa_1_i));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_18 (.A(
        early_flags_pmux_63_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[60]), .D(early_flags_Z[124]), .FCI(
        early_flags_pmux_63_1_1_co0_8), .S(
        early_flags_pmux_63_1_1_wmux_18_S_0), .Y(
        early_flags_pmux_63_1_1_y7_0), .FCO(
        early_flags_pmux_63_1_1_co1_8));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_12 (.A(
        late_flags_pmux_126_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[39]), .D(late_flags_Z[103]), .FCI(
        late_flags_pmux_126_1_0_co0_5), .S(
        late_flags_pmux_126_1_0_wmux_12_S_0), .Y(
        late_flags_pmux_126_1_0_y1_0), .FCO(
        late_flags_pmux_126_1_0_co1_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[105]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[105]), .C(
        un10_early_flags[105]), .Y(late_flags_7_fast_0[105]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_166  (.A(
        late_flags_Z[23]), .B(late_flags_Z[22]), .C(late_flags_Z[21]), 
        .D(late_flags_Z[20]), .Y(calc_done25_166));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[13]), 
        .D(early_flags_Z[77]), .FCI(early_flags_pmux_126_1_1_co1_6), 
        .S(early_flags_pmux_126_1_1_wmux_15_S_0), .Y(
        early_flags_pmux_126_1_1_y0_6), .FCO(
        early_flags_pmux_126_1_1_co0_7));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_177  (.A(
        late_flags_Z[83]), .B(late_flags_Z[82]), .C(late_flags_Z[81]), 
        .D(late_flags_Z[80]), .Y(calc_done25_177));
    CFG4 #( .INIT(16'h4000) )  bitalign_curr_state163 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state163_2), .D(bitalign_curr_state_Z[1]), .Y(
        bitalign_curr_state163_Z));
    CFG3 #( .INIT(8'hFE) )  early_flags_1_sqmuxa_RNIRGCS (.A(
        early_flags_1_sqmuxa_Z), .B(un1_tap_cnt_0_sqmuxa_6_0), .C(
        restart_trng_fg_i), .Y(early_flags_0_sqmuxa_2_i));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_2 (.A(
        late_flags_pmux_126_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[51]), .D(late_flags_Z[115]), .FCI(
        late_flags_pmux_126_1_0_co0_0), .S(
        late_flags_pmux_126_1_0_wmux_2_S_0), .Y(
        late_flags_pmux_126_1_0_0_y3), .FCO(
        late_flags_pmux_126_1_0_co1_0));
    CFG2 #( .INIT(4'h8) )  early_flags_0_sqmuxa (.A(
        bitalign_curr_state153_Z), .B(BIT_ALGN_OOR_0_c), .Y(
        early_flags_0_sqmuxa_Z));
    SLE \late_flags[14]  (.D(late_flags_7_fast_0[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[14]));
    SLE \early_flags[51]  (.D(early_flags_7_fast_0[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[51]));
    SLE \early_flags[10]  (.D(early_flags_7_fast_0[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[10]));
    ARI1 #( .INIT(20'h572D8) )  \tapcnt_final_RNIOTM22[1]  (.A(
        un1_tap_cnt_0_sqmuxa_14_0_0[1]), .B(N_60), .C(tap_cnt_Z[1]), 
        .D(tapcnt_final_Z[1]), .FCI(tap_cnt_17_i_m2_cry_0), .S(N_79), 
        .Y(tapcnt_final_RNIOTM22_Y_0[1]), .FCO(tap_cnt_17_i_m2_cry_1));
    SLE \no_early_no_late_val_st2[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[0]));
    SLE mv_dn_fg (.D(tapcnt_final_upd_3_sqmuxa_1), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(mv_dn_fg_0_sqmuxa_i_0_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(mv_dn_fg_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_72_1 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_1_Z[72]));
    GND GND_Z (.Y(GND));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[11]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[11]), .C(
        un10_early_flags[11]), .Y(early_flags_7_fast_0[11]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_1 (.A(
        un16_tapcnt_final_1), .B(un10_tapcnt_final_1), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_0_Z), .S(
        un16_tapcnt_final_cry_1_S_0), .Y(un16_tapcnt_final_cry_1_Y_0), 
        .FCO(un16_tapcnt_final_cry_1_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_16 (.A(
        late_flags_pmux_126_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[47]), .D(late_flags_Z[111]), .FCI(
        late_flags_pmux_126_1_0_co0_7), .S(
        late_flags_pmux_126_1_0_wmux_16_S_0), .Y(
        late_flags_pmux_126_1_0_y5_0), .FCO(
        late_flags_pmux_126_1_0_co1_7));
    SLE \early_flags[39]  (.D(early_flags_7_fast_0[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[39]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_101 (.A(
        un10_early_flags_1_Z[96]), .B(un10_early_flags_1_Z[5]), .C(
        un10_early_flags_2_0[100]), .Y(un10_early_flags[101]));
    SLE \no_early_no_late_val_st1[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[4]));
    SLE \late_flags[98]  (.D(late_flags_7_fast_0[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[98]));
    SLE \late_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[5])
        );
    SLE \late_flags[44]  (.D(late_flags_7_fast_0[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[44]));
    CFG2 #( .INIT(4'h8) )  un1_retrain_adj_tap (.A(mv_dn_fg_Z), .B(
        mv_up_fg_Z), .Y(un1_retrain_adj_tap_i));
    CFG1 #( .INIT(2'h1) )  \rst_cnt_RNO[0]  (.A(rst_cnt_Z[0]), .Y(
        rst_cnt_s[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[55]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[55]), .C(
        un10_early_flags[55]), .Y(late_flags_7_fast_0[55]));
    SLE \late_flags[105]  (.D(late_flags_7_fast_0[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[105]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_16 (.A(
        late_flags_pmux_63_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[46]), .D(late_flags_Z[110]), .FCI(
        late_flags_pmux_63_1_0_co0_7), .S(
        late_flags_pmux_63_1_0_wmux_16_S_0), .Y(
        late_flags_pmux_63_1_0_y5_0), .FCO(
        late_flags_pmux_63_1_0_co1_7));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_125 (.A(tap_cnt_Z[1]), 
        .B(un10_early_flags_1_Z[5]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[125]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_126_1_1_co1_3), .S(
        late_flags_pmux_126_1_1_wmux_9_S_0), .Y(
        late_flags_pmux_126_1_1_wmux_9_Y_0), .FCO(
        late_flags_pmux_126_1_1_co0_4));
    SLE \early_flags[8]  (.D(early_flags_7_fast_0[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[8]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[89]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[89]), .C(
        un10_early_flags[89]), .Y(late_flags_7_fast_0[89]));
    SLE \late_flags[112]  (.D(late_flags_7_fast_0[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[112]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_40_2_0 (.A(tap_cnt_Z[2]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[40]));
    CFG4 #( .INIT(16'hFD31) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNIEIUK5  (
        .A(rx_trng_done_Z), .B(bitalign_curr_state_Z[2]), .C(
        un1_bitalign_curr_state_14_1_Z), .D(N_83), .Y(N_100));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_44_2_0 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[44]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_12 (.A(
        early_flags_pmux_63_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[38]), .D(early_flags_Z[102]), .FCI(
        early_flags_pmux_63_1_0_co0_5), .S(
        early_flags_pmux_63_1_0_wmux_12_S_0), .Y(
        early_flags_pmux_63_1_0_y1_0), .FCO(
        early_flags_pmux_63_1_0_co1_5));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_24_1 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_1_Z[24]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_4 (.A(
        early_flags_pmux_63_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[40]), .D(early_flags_Z[104]), .FCI(
        early_flags_pmux_63_1_1_co0_1), .S(
        early_flags_pmux_63_1_1_wmux_4_S_0), .Y(
        early_flags_pmux_63_1_1_y5), .FCO(
        early_flags_pmux_63_1_1_co1_1));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[15]), 
        .D(early_flags_Z[79]), .FCI(early_flags_pmux_126_1_0_co1_6), 
        .S(early_flags_pmux_126_1_0_wmux_15_S_0), .Y(
        early_flags_pmux_126_1_0_y0_6), .FCO(
        early_flags_pmux_126_1_0_co0_7));
    SLE \early_flags[84]  (.D(early_flags_7_fast_0[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[84]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_136  (.A(
        early_flags_Z[87]), .B(early_flags_Z[86]), .C(
        early_flags_Z[85]), .D(early_flags_Z[84]), .Y(calc_done25_136));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[4]), 
        .D(early_flags_Z[68]), .FCI(early_flags_pmux_63_1_1_co1_4), .S(
        early_flags_pmux_63_1_1_wmux_11_S_0), .Y(
        early_flags_pmux_63_1_1_y0_4), .FCO(
        early_flags_pmux_63_1_1_co0_5));
    CFG4 #( .INIT(16'hFE00) )  bitalign_curr_state12_0_0 (.A(
        BIT_ALGN_EYE_IN_c[2]), .B(BIT_ALGN_EYE_IN_c[1]), .C(
        BIT_ALGN_EYE_IN_c[0]), .D(PLL_LOCK_0), .Y(
        bitalign_curr_state12_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[26]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[26]), .C(
        un10_early_flags[26]), .Y(early_flags_7_fast_0[26]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_28_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[1]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[28]));
    CFG4 #( .INIT(16'hF5F4) )  \un1_tap_cnt_0_sqmuxa_14_0[1]  (.A(
        un1_early_flags_1_sqmuxa_i), .B(N_82), .C(restart_trng_fg_i), 
        .D(bitalign_curr_state_0_sqmuxa_10), .Y(
        un1_tap_cnt_0_sqmuxa_14_0_0[1]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[86]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[86]), .C(
        un10_early_flags[86]), .Y(early_flags_7_fast_0[86]));
    SLE \early_flags[69]  (.D(early_flags_7_fast_0[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[69]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[93]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[93]), .C(
        un10_early_flags[93]), .Y(late_flags_7_fast_0[93]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI3CJ81[2]  (.A(early_val_Z[2])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[2]), .Y(
        early_val_RNI3CJ81_Z[2]));
    SLE \early_flags[12]  (.D(early_flags_7_fast_0[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[12]));
    CFG4 #( .INIT(16'hDFFF) )  \late_flags_7_i_o4[49]  (.A(
        tap_cnt_Z[0]), .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[48]), 
        .D(un10_early_flags_1_Z[48]), .Y(N_208));
    SLE \no_early_no_late_val_st2[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[3]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_101_2 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[6]), .Y(un10_early_flags_1_Z[96]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[26]), 
        .D(late_flags_Z[90]), .FCI(late_flags_pmux_63_1_0_co1_1), .S(
        late_flags_pmux_63_1_0_wmux_5_S_0), .Y(
        late_flags_pmux_63_1_0_y0_2), .FCO(
        late_flags_pmux_63_1_0_co0_2));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_48_1 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[4]), .Y(un10_early_flags_1_Z[48]));
    CFG2 #( .INIT(4'h7) )  un10_early_flags_18_1_i (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[1]), .Y(N_1499));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[120]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[120]), .C(
        un10_early_flags[120]), .Y(late_flags_7_fast_0[120]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_7 (.A(
        early_flags_pmux_63_1_0_0_y7), .B(early_flags_pmux_63_1_0_0_y5)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co1_2), .S(
        early_flags_pmux_63_1_0_wmux_7_S_0), .Y(
        early_flags_pmux_63_1_0_y0_3), .FCO(
        early_flags_pmux_63_1_0_co0_3));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_92 (.A(
        un10_early_flags_1_Z[12]), .B(un10_early_flags_1_Z[0]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_1_Z[80]), .Y(
        un10_early_flags[92]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[66]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[66]), .C(
        un10_early_flags[66]), .Y(early_flags_7_fast_0[66]));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_start_7_s_7 (.A(
        VCC), .B(un1_restart_trng_fg_5_0), .C(GND), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_6), .S(
        noearly_nolate_diff_start_7[7]), .Y(
        noearly_nolate_diff_start_7_s_7_Y_0), .FCO(
        noearly_nolate_diff_start_7_s_7_FCO_0));
    CFG2 #( .INIT(4'h8) )  tap_cnt_0_sqmuxa_1 (.A(
        bitalign_curr_state148_Z), .B(bitalign_curr_state12_Z), .Y(
        tap_cnt_0_sqmuxa_1_Z));
    SLE mv_up_fg (.D(tapcnt_final_upd_2_sqmuxa_1), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(mv_up_fg_0_sqmuxa_i_0_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(mv_up_fg_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_164  (.A(
        late_flags_Z[31]), .B(late_flags_Z[30]), .C(late_flags_Z[29]), 
        .D(late_flags_Z[28]), .Y(calc_done25_164));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_74 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_1_Z[10]), .C(
        un10_early_flags_2_0[72]), .Y(un10_early_flags[74]));
    SLE \late_flags[2]  (.D(late_flags_7_fast_0[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[2]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI9ABM[0]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[0]), .D(GND), .FCI(
        timeout_cnt_cry_cy), .S(timeout_cnt_s[0]), .Y(
        timeout_cnt_RNI9ABM_Y_0[0]), .FCO(timeout_cnt_cry[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_4 (.A(
        late_flags_pmux_126_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[41]), .D(late_flags_Z[105]), .FCI(
        late_flags_pmux_126_1_1_co0_1), .S(
        late_flags_pmux_126_1_1_wmux_4_S_0), .Y(
        late_flags_pmux_126_1_1_y5), .FCO(
        late_flags_pmux_126_1_1_co1_1));
    SLE \early_flags[86]  (.D(early_flags_7_fast_0[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[86]));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_start_7_cry_0_0_cy 
        (.A(VCC), .B(un1_restart_trng_fg_5_0), .C(GND), .D(GND), .FCI(
        VCC), .S(noearly_nolate_diff_start_7_cry_0_0_cy_S_0), .Y(
        noearly_nolate_diff_start_7_cry_0_0_cy_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_0_0_cy_Z));
    SLE \early_flags[9]  (.D(early_flags_7_fast_0[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[9]));
    SLE \early_flags[94]  (.D(early_flags_7_fast_0[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[94]));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_113 (.A(tap_cnt_Z[3]), 
        .B(N_1498), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[113]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[75]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[75]), .C(
        un10_early_flags[75]), .Y(late_flags_7_fast_0[75]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[86]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[86]), .C(
        un10_early_flags[86]), .Y(late_flags_7_fast_0[86]));
    SLE \early_flags[87]  (.D(early_flags_7_fast_0[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[87]));
    SLE \late_flags[127]  (.D(late_flags_7_fast_0[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[127]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_10 (.A(
        late_flags_pmux_63_1_1_y21), .B(late_flags_pmux_63_1_1_y9), .C(
        emflag_cnt_Z[2]), .D(VCC), .FCI(late_flags_pmux_63_1_1_co0_4), 
        .S(late_flags_pmux_63_1_1_wmux_10_S_0), .Y(
        late_flags_pmux_63_1_1_wmux_10_Y_0), .FCO(
        late_flags_pmux_63_1_1_co1_4));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[125]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[125]), .C(
        un10_early_flags[125]), .Y(late_flags_7_fast_0[125]));
    SLE rx_trng_done (.D(N_1403), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(rx_trng_done_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_trng_done_Z));
    SLE \late_flags[94]  (.D(late_flags_7_fast_0[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[94]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[68]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[68]), .C(
        un10_early_flags[68]), .Y(late_flags_7_fast_0[68]));
    CFG3 #( .INIT(8'hC8) )  
        \bitalign_curr_state_34_4_0_.un1_bitalign_curr_state_2_sqmuxa  
        (.A(emflag_cnt_0_sqmuxa), .B(bitalign_curr_state89), .C(
        bitalign_curr_state159), .Y(un1_bitalign_curr_state_2_sqmuxa));
    SLE \early_flags[81]  (.D(early_flags_7_fast_0[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[81]));
    SLE late_cur_set (.D(late_cur_set_2_sqmuxa), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(late_cur_set_0_sqmuxa_i), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(late_cur_set_Z));
    SLE \early_flags[79]  (.D(early_flags_7_fast_0[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[79]));
    CFG4 #( .INIT(16'hFFFE) )  bitalign_curr_state61_NE_4 (.A(
        bitalign_curr_state61_6_Z), .B(bitalign_curr_state61_3_Z), .C(
        bitalign_curr_state61_2_Z), .D(bitalign_curr_state61_1_Z), .Y(
        bitalign_curr_state61_NE_4_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[106]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[106]), .C(
        un10_early_flags[106]), .Y(early_flags_7_fast_0[106]));
    SLE \retrain_reg[2]  (.D(retrain_reg_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(retrain_reg_Z[2]));
    CFG2 #( .INIT(4'hD) )  \bitalign_curr_state_34_4_0_.m68  (.A(
        bitalign_curr_state13), .B(bitalign_curr_state_Z[0]), .Y(N_69));
    SLE \late_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[1])
        );
    CFG2 #( .INIT(4'h1) )  un10_early_flags_0_1 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_1_Z[0]));
    CFG3 #( .INIT(8'h10) )  mv_dn_fg_0_sqmuxa_i_a2_0_RNIHVRK (.A(
        mv_up_fg_Z), .B(bitalign_curr_state12_Z), .C(N_98), .Y(
        tapcnt_final_upd_1_sqmuxa));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[112]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[112]), .C(
        un10_early_flags[112]), .Y(early_flags_7_fast_0[112]));
    SLE \early_flags[104]  (.D(early_flags_7_fast_0[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[104]));
    SLE \emflag_cnt[3]  (.D(emflag_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[58]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[58]), .C(
        un10_early_flags[58]), .Y(early_flags_7_fast_0[58]));
    ARI1 #( .INIT(20'h51144) )  tapcnt_final_upd_8_cry_2_0 (.A(
        tapcnt_final_upd_1_sqmuxa), .B(mv_dn_fg_0_sqmuxa_i_o2_0), .C(
        tap_cnt_Z[2]), .D(GND), .FCI(GND), .S(
        tapcnt_final_upd_8_cry_2_0_S_0), .Y(
        tapcnt_final_upd_8_cry_2_0_Y_0), .FCO(tapcnt_final_upd_8_cry_2)
        );
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[1]  (.A(VCC), .B(
        rst_cnt_Z[1]), .C(GND), .D(GND), .FCI(rst_cnt_s_715_FCO_0), .S(
        rst_cnt_s[1]), .Y(rst_cnt_cry_Y_1[1]), .FCO(rst_cnt_cry_Z[1]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_21_2 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[21]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_80_1 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[4]), .Y(un10_early_flags_1_Z[80]));
    SLE \no_early_no_late_val_end1[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[57]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[57]), .C(
        un10_early_flags[57]), .Y(late_flags_7_fast_0[57]));
    ARI1 #( .INIT(20'h45500) )  early_late_diff_8_s_7 (.A(VCC), .B(
        un1_restart_trng_fg_5_0), .C(GND), .D(GND), .FCI(
        early_late_diff_8_cry_6), .S(early_late_diff_8[7]), .Y(
        early_late_diff_8_s_7_Y_0), .FCO(early_late_diff_8_s_7_FCO_0));
    SLE \tapcnt_final_upd[5]  (.D(tapcnt_final_upd_8[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[5]));
    SLE \noearly_nolate_diff_start[5]  (.D(
        noearly_nolate_diff_start_7[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_5));
    SLE \early_flags[58]  (.D(early_flags_7_fast_0[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[58]));
    CFG4 #( .INIT(16'h1300) )  \bitalign_curr_state_34_4_0_.m19  (.A(
        late_cur_set_Z), .B(early_cur_set_Z), .C(late_flags_pmux), .D(
        early_flags_pmux), .Y(N_20));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[55]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[55]), .C(
        un10_early_flags[55]), .Y(early_flags_7_fast_0[55]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_134  (.A(
        early_flags_Z[111]), .B(early_flags_Z[110]), .C(
        early_flags_Z[109]), .D(early_flags_Z[108]), .Y(
        calc_done25_134));
    SLE \early_flags[96]  (.D(early_flags_7_fast_0[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[96]));
    SLE \emflag_cnt[2]  (.D(emflag_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[5]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[5]), .C(
        un10_early_flags[5]), .Y(early_flags_7_fast_0[5]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[16]), 
        .D(late_flags_Z[80]), .FCI(late_flags_pmux_63_1_1_co1), .S(
        late_flags_pmux_63_1_1_wmux_1_S_0), .Y(
        late_flags_pmux_63_1_1_y0_0), .FCO(
        late_flags_pmux_63_1_1_co0_0));
    SLE \early_flags[97]  (.D(early_flags_7_fast_0[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[97]));
    SLE \early_flags[126]  (.D(early_flags_7_fast_0[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[126]));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_4 (.A(
        tapcnt_final_upd_Z[4]), .B(tapcnt_final_Z[4]), .C(tap_cnt_Z[4])
        , .D(N_1416), .Y(bitalign_curr_state61_4_Z));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_64_1 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[64]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[101]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[101]), .C(
        un10_early_flags[101]), .Y(late_flags_7_fast_0[101]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_103 (.A(
        un10_early_flags_1_Z[36]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_3_Z[87]), .Y(
        un10_early_flags[103]));
    CFG3 #( .INIT(8'h27) )  \bitalign_curr_state_34_4_0_.m23_1_2  (.A(
        late_last_set15_Z), .B(late_flags_pmux), .C(N_20), .Y(m23_1_2));
    CFG4 #( .INIT(16'h2000) )  bitalign_curr_state162 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state161_2_Z), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state162_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[105]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[105]), .C(
        un10_early_flags[105]), .Y(early_flags_7_fast_0[105]));
    SLE \late_flags[5]  (.D(late_flags_7_fast_0[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[104]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[104]), .C(
        un10_early_flags[104]), .Y(early_flags_7_fast_0[104]));
    SLE \early_flags[91]  (.D(early_flags_7_fast_0[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[91]));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[4]  (.A(
        tapcnt_final_13_Z[5]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[4]), .Y(tapcnt_final_13_1_Z[4]));
    SLE \late_flags[26]  (.D(late_flags_7_fast_0[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[26]));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[4]  (.A(
        no_early_no_late_val_end1_Z[4]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[4]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[4]));
    ARI1 #( .INIT(20'h54411) )  tapcnt_final_upd_8_cry_3_0 (.A(
        tap_cnt_Z[3]), .B(mv_dn_fg_0_sqmuxa_i_o2_0), .C(
        tapcnt_final_upd_1_sqmuxa), .D(GND), .FCI(
        tapcnt_final_upd_8_cry_2), .S(tapcnt_final_upd_8[3]), .Y(
        tapcnt_final_upd_8_cry_3_0_Y_0), .FCO(tapcnt_final_upd_8_cry_3)
        );
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[48]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[48]), .C(
        un10_early_flags[48]), .Y(early_flags_7_fast_0[48]));
    CFG4 #( .INIT(16'hCCEC) )  un1_tap_cnt_0_sqmuxa_1 (.A(
        bitalign_curr_state149_Z), .B(tap_cnt_0_sqmuxa_1_Z), .C(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .D(BIT_ALGN_ERR_c), .Y(
        un1_tap_cnt_0_sqmuxa_6_0));
    CFG3 #( .INIT(8'h80) )  \bitalign_curr_state_34_4_0_.calc_done25  
        (.A(calc_done25_248), .B(calc_done25_253), .C(calc_done25_249), 
        .Y(calc_done25));
    CFG4 #( .INIT(16'h71F9) )  \bitalign_curr_state_34_4_0_.m37_1_1  (
        .A(bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[0]), .C(
        early_flags_pmux), .D(N_35), .Y(m37_1_1));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_3 (.A(
        un16_tapcnt_final_3), .B(un10_tapcnt_final_3), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_2_Z), .S(
        un16_tapcnt_final_cry_3_S_0), .Y(un16_tapcnt_final_cry_3_Y_0), 
        .FCO(un16_tapcnt_final_cry_3_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_43 (.A(
        un10_early_flags_2_0[40]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[40]), .Y(un10_early_flags[43]));
    SLE \wait_cnt[1]  (.D(wait_cnt_4_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(wait_cnt_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[99]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[99]), .C(
        un10_early_flags[99]), .Y(late_flags_7_fast_0[99]));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[5]  (.A(
        tapcnt_final_13_Z[6]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[5]), .Y(tapcnt_final_13_1_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[45]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[45]), .C(
        un10_early_flags[45]), .Y(early_flags_7_fast_0[45]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_89 (.A(tap_cnt_Z[5]), 
        .B(un10_early_flags_1_Z[9]), .C(un10_early_flags_1_Z[80]), .D(
        un10_early_flags_2_Z[8]), .Y(un10_early_flags[89]));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_nxt_8_s_7 (.A(VCC), 
        .B(un1_restart_trng_fg_5_0), .C(GND), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_6), .S(
        noearly_nolate_diff_nxt_8[7]), .Y(
        noearly_nolate_diff_nxt_8_s_7_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_s_7_FCO_0));
    CFG4 #( .INIT(16'hFEFF) )  un1_bitalign_curr_state_12 (.A(
        early_flags_1_sqmuxa_1_Z), .B(early_flags_0_sqmuxa_1_Z), .C(
        bitalign_curr_state_Z[1]), .D(un1_bitalign_curr_state148_3_Z), 
        .Y(un1_bitalign_curr_state_12_Z));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state_0_sqmuxa_9 (.A(
        rx_err_1_sqmuxa_Z), .B(calc_done_4_sqmuxa_0_Z), .C(
        un1_bitalign_curr_state_0_sqmuxa_9_4_Z), .Y(
        un1_bitalign_curr_state_0_sqmuxa_9_i));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[118]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[118]), .C(
        un10_early_flags[118]), .Y(early_flags_7_fast_0[118]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_181  (.A(
        late_flags_Z[75]), .B(late_flags_Z[74]), .C(late_flags_Z[73]), 
        .D(late_flags_Z[72]), .Y(calc_done25_181));
    CFG4 #( .INIT(16'h1000) )  bitalign_curr_state156 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state152_1_Z), .D(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state156_Z));
    CFG4 #( .INIT(16'h0080) )  bitalign_curr_state_0_sqmuxa_8 (.A(
        bitalign_curr_state41_Z), .B(bitalign_curr_state152_3_Z), .C(
        BIT_ALGN_OOR_0_c), .D(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state_0_sqmuxa_8_Z));
    SLE \late_flags[76]  (.D(late_flags_7_fast_0[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[76]));
    CFG2 #( .INIT(4'h2) )  \bitalign_curr_state_34_4_0_.m55_0  (.A(
        bitalign_curr_state161_2_Z), .B(bitalign_curr_state_Z[0]), .Y(
        m55_0));
    CFG2 #( .INIT(4'h2) )  early_late_diff_2_sqmuxa (.A(
        early_late_diff_0_sqmuxa_Z), .B(restart_trng_fg_i), .Y(
        early_late_diff_2_sqmuxa_Z));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_95 (.A(
        un10_early_flags_1_Z[80]), .B(tap_cnt_Z[5]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[95]));
    CFG3 #( .INIT(8'h10) )  \bitalign_curr_state_34_4_0_.m52  (.A(
        late_last_set15_Z), .B(early_flags_dec[127]), .C(N_20), .Y(
        N_119_mux));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[77]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[77]), .C(
        un10_early_flags[77]), .Y(late_flags_7_fast_0[77]));
    CFG4 #( .INIT(16'h00CA) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNIBD2F5  (
        .A(i22_mux), .B(N_130_mux), .C(bitalign_curr_state_Z[4]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[4]));
    SLE reset_dly_fg (.D(VCC), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(reset_dly_fg4_Z), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(reset_dly_fg_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_0 (.A(
        late_flags_pmux_63_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[32]), .D(late_flags_Z[96]), .FCI(
        late_flags_pmux_63_1_1_co0), .S(
        late_flags_pmux_63_1_1_wmux_0_S_0), .Y(
        late_flags_pmux_63_1_1_y1), .FCO(late_flags_pmux_63_1_1_co1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[111]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[111]), .C(
        un10_early_flags[111]), .Y(early_flags_7_fast_0[111]));
    ARI1 #( .INIT(20'h0FA44) )  
        \bitalign_curr_state_34_4_0_.m74_2_1_1_1_wmux  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        N_69), .D(m74_1_0_0), .FCI(VCC), .S(m74_2_1_1_wmux_S_0), .Y(
        m74_2_1_1_1_y0), .FCO(m74_2_1_1_1_co0));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_8_2 (.A(tap_cnt_Z[1]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[8]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[32]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[32]), .C(
        un10_early_flags[32]), .Y(early_flags_7_fast_0[32]));
    CFG4 #( .INIT(16'hFFFE) )  un2_early_late_diff_validlto7_2 (.A(
        early_late_diff_Z[7]), .B(early_late_diff_Z[6]), .C(
        early_late_diff_Z[5]), .D(early_late_diff_Z[4]), .Y(
        un2_early_late_diff_validlto7_2_Z));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_1_wmux_8 (.A(
        late_flags_pmux_126_1_1_y0_3), .B(late_flags_pmux_126_1_1_y3), 
        .C(late_flags_pmux_126_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co0_3), .S(
        late_flags_pmux_126_1_1_wmux_8_S_0), .Y(
        late_flags_pmux_126_1_1_y9), .FCO(
        late_flags_pmux_126_1_1_co1_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[31]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[31]), .C(
        un10_early_flags[31]), .Y(late_flags_7_fast_0[31]));
    SLE \late_flags[7]  (.D(late_flags_7_fast_0[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[7]));
    CFG4 #( .INIT(16'h0400) )  \bitalign_curr_state_34_4_0_.m91_2  (.A(
        bitalign_curr_state_Z[1]), .B(tap_cnt_0_sqmuxa_0_Z), .C(
        calc_done_Z), .D(bitalign_curr_state_Z[2]), .Y(m91_1));
    SLE \late_flags[36]  (.D(late_flags_7_fast_0[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[36]));
    SLE \late_flags[57]  (.D(late_flags_7_fast_0[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[57]));
    CFG4 #( .INIT(16'hF2F0) )  un1_early_flags_1_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(mv_dn_fg_Z), .C(
        early_flags_1_sqmuxa_Z), .D(bitalign_curr_state156_Z), .Y(
        un1_early_flags_1_sqmuxa_i));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_32 (.A(
        un10_early_flags_1_Z[32]), .B(un10_early_flags_2_Z[8]), .C(
        un10_early_flags_2_0[32]), .Y(un10_early_flags[32]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[11]), 
        .D(late_flags_Z[75]), .FCI(late_flags_pmux_126_1_0_co1_0), .S(
        late_flags_pmux_126_1_0_wmux_3_S_0), .Y(
        late_flags_pmux_126_1_0_y0_1), .FCO(
        late_flags_pmux_126_1_0_co0_1));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_5_0 (.A(
        emflag_cnt_Z[5]), .B(un1_restart_trng_fg_5_0), .C(
        early_val_Z[5]), .D(GND), .FCI(early_late_diff_8_cry_4), .S(
        early_late_diff_8[5]), .Y(early_late_diff_8_cry_5_0_Y_0), .FCO(
        early_late_diff_8_cry_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[21]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[21]), .C(
        un10_early_flags[21]), .Y(late_flags_7_fast_0[21]));
    SLE \late_flags[21]  (.D(late_flags_7_fast_0[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[21]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[1]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[1]), .D(GND), .FCI(
        emflag_cnt_cry_Z[0]), .S(emflag_cnt_s[1]), .Y(
        emflag_cnt_cry_Y_1[1]), .FCO(emflag_cnt_cry_Z[1]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_3 (.A(
        un10_tapcnt_final_3), .B(early_late_diff_Z[3]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_2_Z), .S(
        un1_early_late_diff_cry_3_S_0), .Y(
        un1_early_late_diff_cry_3_Y_0), .FCO(
        un1_early_late_diff_cry_3_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[96]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[96]), .C(
        un10_early_flags[96]), .Y(late_flags_7_fast_0[96]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[1]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[1]), .C(
        un10_early_flags[1]), .Y(late_flags_7_fast_0[1]));
    CFG4 #( .INIT(16'h0008) )  bit_align_dly_done_0_sqmuxa_1_0 (.A(
        rx_trng_done_Z), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state_Z[4]), .D(bitalign_curr_state_Z[0]), .Y(
        bit_align_dly_done_0_sqmuxa_1_0_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[96]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[96]), .C(
        un10_early_flags[96]), .Y(early_flags_7_fast_0[96]));
    SLE \tapcnt_final[6]  (.D(tapcnt_final_13_1_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[0]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[0]), .C(
        un10_early_flags[0]), .Y(late_flags_7_fast_0[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_14 (.A(
        late_flags_pmux_126_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[53]), .D(late_flags_Z[117]), .FCI(
        late_flags_pmux_126_1_1_co0_6), .S(
        late_flags_pmux_126_1_1_wmux_14_S_0), .Y(
        late_flags_pmux_126_1_1_y3_0), .FCO(
        late_flags_pmux_126_1_1_co1_6));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_77 (.A(
        un10_early_flags_2_0[76]), .B(un10_early_flags_1_Z[72]), .C(
        un10_early_flags_1_Z[5]), .Y(un10_early_flags[77]));
    CFG4 #( .INIT(16'hF400) )  bit_align_done_0_sqmuxa_2 (.A(
        un1_retrain_adj_tap_i), .B(un1_rx_BIT_ALGN_START), .C(
        bitalign_curr_state12_Z), .D(bitalign_curr_state148_Z), .Y(
        bit_align_done_0_sqmuxa_2_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[17]), 
        .D(late_flags_Z[81]), .FCI(late_flags_pmux_126_1_1_co1), .S(
        late_flags_pmux_126_1_1_wmux_1_S_0), .Y(
        late_flags_pmux_126_1_1_y0_0), .FCO(
        late_flags_pmux_126_1_1_co0_0));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_3 (.A(
        tapcnt_final_upd_Z[3]), .B(tapcnt_final_Z[3]), .C(tap_cnt_Z[3])
        , .D(N_1416), .Y(bitalign_curr_state61_3_Z));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI8UO41[1]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[1]), .D(GND), .FCI(
        timeout_cnt_cry[0]), .S(timeout_cnt_s[1]), .Y(
        timeout_cnt_RNI8UO41_Y_0[1]), .FCO(timeout_cnt_cry[1]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_96_2_0 (.A(
        un10_early_flags_2_Z[0]), .B(tap_cnt_Z[4]), .Y(
        un10_early_flags_2_0[96]));
    SLE \early_flags[88]  (.D(early_flags_7_fast_0[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[88]));
    SLE \early_late_diff[0]  (.D(early_late_diff_8[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[0]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_0 (.A(
        un10_tapcnt_final_0), .B(un16_tapcnt_final_0), .C(GND), .D(GND)
        , .FCI(GND), .S(un10_tapcnt_final_cry_0_S_0), .Y(
        un10_tapcnt_final_cry_0_Y_0), .FCO(un10_tapcnt_final_cry_0_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_167  (.A(
        late_flags_Z[19]), .B(late_flags_Z[18]), .C(late_flags_Z[17]), 
        .D(late_flags_Z[16]), .Y(calc_done25_167));
    SLE \noearly_nolate_diff_nxt[6]  (.D(noearly_nolate_diff_nxt_8[6]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_6));
    CFG4 #( .INIT(16'h0002) )  \tapcnt_final_13_sn.m6  (.A(
        calc_done_4_sqmuxa_0_Z), .B(un1_calc_done25_5), .C(
        tapcnt_final27), .D(restart_trng_fg_i), .Y(
        tapcnt_final_5_sqmuxa));
    SLE \tapcnt_final[1]  (.D(tapcnt_final_13_1_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[1]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_0 (.A(
        late_flags_pmux_126_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[35]), .D(late_flags_Z[99]), .FCI(
        late_flags_pmux_126_1_0_0_co0), .S(
        late_flags_pmux_126_1_0_wmux_0_S_0), .Y(
        late_flags_pmux_126_1_0_0_y1), .FCO(
        late_flags_pmux_126_1_0_0_co1));
    SLE \cnt[1]  (.D(cnt_RNO_0[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(cnt_Z[1]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_22 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_2_0[16]), .C(
        un10_early_flags_1_Z[16]), .Y(un10_early_flags[22]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[121]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[121]), .C(
        un10_early_flags[121]), .Y(late_flags_7_fast_0[121]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[9]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[9]), .C(
        un10_early_flags[9]), .Y(late_flags_7_fast_0[9]));
    SLE \late_flags[4]  (.D(late_flags_7_fast_0[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[4]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_0_0 (
        .A(emflag_cnt_Z[0]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st1_Z[0]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_0_0_cy_Z), .S(
        noearly_nolate_diff_start_7[0]), .Y(
        noearly_nolate_diff_start_7_cry_0_0_Y_0), .FCO(
        noearly_nolate_diff_start_7_cry_0));
    SLE \late_flags[71]  (.D(late_flags_7_fast_0[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[71]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[7]), 
        .D(early_flags_Z[71]), .FCI(early_flags_pmux_126_1_0_co1_4), 
        .S(early_flags_pmux_126_1_0_wmux_11_S_0), .Y(
        early_flags_pmux_126_1_0_y0_4), .FCO(
        early_flags_pmux_126_1_0_co0_5));
    CFG4 #( .INIT(16'h4073) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNISBQ9B  (
        .A(bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        N_100), .D(m101_1_1), .Y(N_102));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_2 (.A(
        early_flags_pmux_63_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[50]), .D(early_flags_Z[114]), .FCI(
        early_flags_pmux_63_1_0_co0_0), .S(
        early_flags_pmux_63_1_0_wmux_2_S_0), .Y(
        early_flags_pmux_63_1_0_0_y3), .FCO(
        early_flags_pmux_63_1_0_co1_0));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[27]), 
        .D(early_flags_Z[91]), .FCI(early_flags_pmux_126_1_0_co1_1), 
        .S(early_flags_pmux_126_1_0_wmux_5_S_0), .Y(
        early_flags_pmux_126_1_0_y0_2), .FCO(
        early_flags_pmux_126_1_0_co0_2));
    SLE \early_flags[1]  (.D(early_flags_7_fast_0[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[1]));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_0_2 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[53]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[53]), .C(
        un10_early_flags[53]), .Y(early_flags_7_fast_0[53]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[41]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[41]), .C(
        un10_early_flags[41]), .Y(late_flags_7_fast_0[41]));
    SLE \tapcnt_final[5]  (.D(tapcnt_final_13_1_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[27]), 
        .D(late_flags_Z[91]), .FCI(late_flags_pmux_126_1_0_co1_1), .S(
        late_flags_pmux_126_1_0_wmux_5_S_0), .Y(
        late_flags_pmux_126_1_0_y0_2), .FCO(
        late_flags_pmux_126_1_0_co0_2));
    SLE \late_flags[67]  (.D(late_flags_7_fast_0[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[67]));
    SLE \no_early_no_late_val_end2[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[4]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_98 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_1_Z[64]), .D(
        un10_early_flags_2_0[96]), .Y(un10_early_flags[98]));
    CFG3 #( .INIT(8'hEA) )  un2_noearly_nolate_diff_nxt_validlto2 (.A(
        un16_tapcnt_final_2), .B(un16_tapcnt_final_1), .C(
        un16_tapcnt_final_0), .Y(un2_noearly_nolate_diff_nxt_validlt3));
    SLE \restart_reg[0]  (.D(debouncer_0_DB_OUT), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_reg_Z[0]));
    SLE \early_flags[35]  (.D(early_flags_7_fast_0[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[35]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_19 (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[16]), .Y(un10_early_flags[19]));
    CFG4 #( .INIT(16'hCA42) )  \bitalign_curr_state_34_4_0_.m64  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        m64_1_1), .D(N_63), .Y(N_65));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_5 (.A(
        un16_tapcnt_final_5), .B(early_late_diff_Z[5]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_4_Z), .S(
        un1_early_late_diff_1_cry_5_S_0), .Y(
        un1_early_late_diff_1_cry_5_Y_0), .FCO(
        un1_early_late_diff_1_cry_5_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_9 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_126_1_1_co1_3), .S(
        early_flags_pmux_126_1_1_wmux_9_S_0), .Y(
        early_flags_pmux_126_1_1_wmux_9_Y_0), .FCO(
        early_flags_pmux_126_1_1_co0_4));
    SLE \late_flags[80]  (.D(late_flags_7_fast_0[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[80]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_156  (.A(
        early_flags_Z[15]), .B(early_flags_Z[14]), .C(
        early_flags_Z[13]), .D(early_flags_Z[12]), .Y(calc_done25_156));
    CFG2 #( .INIT(4'h2) )  bit_align_dly_done_2_sqmuxa (.A(
        bitalign_curr_state_0_sqmuxa_9_Z), .B(restart_trng_fg_i), .Y(
        bit_align_dly_done_2_sqmuxa_Z));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_183  (.A(
        late_flags_Z[71]), .B(late_flags_Z[70]), .C(late_flags_Z[69]), 
        .D(late_flags_Z[68]), .Y(calc_done25_183));
    CFG2 #( .INIT(4'hE) )  un1_bitalign_curr_state148_8_1 (.A(
        early_flags_1_sqmuxa_1_Z), .B(early_flags_0_sqmuxa_1_Z), .Y(
        un1_bitalign_curr_state148_8_1_Z));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIRRPT[4]  (.A(
        no_early_no_late_val_st1_Z[4]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_st2_Z[4]), .Y(
        un1_no_early_no_late_val_st1_1_1[4]));
    SLE \late_flags[31]  (.D(late_flags_7_fast_0[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[31]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[117]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[117]), .C(
        un10_early_flags[117]), .Y(early_flags_7_fast_0[117]));
    SLE \early_flags[98]  (.D(early_flags_7_fast_0[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[98]));
    CFG4 #( .INIT(16'h0421) )  un1_bitalign_curr_state148_3 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state_Z[0]), .D(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state148_3_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_76 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_2_0[76]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[76]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_239  (.A(
        calc_done25_191), .B(calc_done25_190), .C(calc_done25_189), .D(
        calc_done25_188), .Y(calc_done25_239));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_115 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_2_Z[67]), .Y(
        un10_early_flags[115]));
    SLE \no_early_no_late_val_st1[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[0]));
    CFG4 #( .INIT(16'hFFF1) )  un1_bitalign_curr_state148_8_2 (.A(
        un1_bitalign_curr_state148_5_4_Z), .B(
        un1_bitalign_curr_state148_4_1_Z), .C(
        un1_bitalign_curr_state148_8_0_Z), .D(rx_trng_done_1_sqmuxa_Z), 
        .Y(un1_bitalign_curr_state148_8_2_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_4 (.A(
        late_flags_pmux_63_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[42]), .D(late_flags_Z[106]), .FCI(
        late_flags_pmux_63_1_0_co0_1), .S(
        late_flags_pmux_63_1_0_wmux_4_S_0), .Y(
        late_flags_pmux_63_1_0_0_y5), .FCO(
        late_flags_pmux_63_1_0_co1_1));
    CFG4 #( .INIT(16'h0080) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state89_RNIQCDC5  (
        .A(bitalign_curr_state_Z[2]), .B(N_83), .C(
        bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[4]), .Y(
        m85_1));
    SLE \rst_cnt[5]  (.D(rst_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[5]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_137  (.A(
        early_flags_Z[83]), .B(early_flags_Z[82]), .C(
        early_flags_Z[81]), .D(early_flags_Z[80]), .Y(calc_done25_137));
    CFG4 #( .INIT(16'hFF8C) )  un1_restart_trng_fg_10 (.A(calc_done25), 
        .B(bitalign_curr_state162_Z), .C(un1_calc_done25_7_i), .D(
        un1_restart_trng_fg_10_0_Z), .Y(un1_restart_trng_fg_10_sn));
    SLE \tap_cnt[0]  (.D(N_32_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[0]));
    SLE \no_early_no_late_val_end1[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[33]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[33]), .C(
        un10_early_flags[33]), .Y(late_flags_7_fast_0[33]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[43]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[43]), .C(
        un10_early_flags[43]), .Y(early_flags_7_fast_0[43]));
    SLE \late_flags[10]  (.D(late_flags_7_fast_0[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[10]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_190  (.A(
        late_flags_Z[111]), .B(late_flags_Z[110]), .C(
        late_flags_Z[109]), .D(late_flags_Z[108]), .Y(calc_done25_190));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[102]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[102]), .C(
        un10_early_flags[102]), .Y(early_flags_7_fast_0[102]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_7 (.A(
        un10_tapcnt_final_7), .B(un16_tapcnt_final_7), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_6_Z), .S(
        un10_tapcnt_final_cry_7_S_0), .Y(un10_tapcnt_final_cry_7_Y_0), 
        .FCO(un10_tapcnt_final_cry_7_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_6_1 (.A(tap_cnt_Z[1]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[6]));
    SLE \early_flags[65]  (.D(early_flags_7_fast_0[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[65]));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[3]  (.A(N_77), .B(N_63_0), .Y(
        N_26_i));
    ARI1 #( .INIT(20'h572D8) )  \tapcnt_final_RNI2SF33[2]  (.A(
        un1_tap_cnt_0_sqmuxa_14_0_0[1]), .B(N_60), .C(tap_cnt_Z[2]), 
        .D(tapcnt_final_Z[2]), .FCI(tap_cnt_17_i_m2_cry_1), .S(N_78), 
        .Y(tapcnt_final_RNI2SF33_Y_0[2]), .FCO(tap_cnt_17_i_m2_cry_2));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNISIPVK[5]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIROIR_0[5]), .B(
        early_val_RNICLJ81_Z[5]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[5]), .FCI(tapcnt_final_13_m1_cry_4), .S(
        tapcnt_final_13_m1[5]), .Y(early_val_RNISIPVK_Y[5]), .FCO(
        tapcnt_final_13_m1_cry_5));
    SLE \bitalign_curr_state[2]  (.D(bitalign_curr_state_34[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[2]));
    ARI1 #( .INIT(20'h574B8) )  \tapcnt_final_RNIES844[3]  (.A(
        tap_cnt_Z[3]), .B(un1_tap_cnt_0_sqmuxa_14_0_0[1]), .C(N_60), 
        .D(tapcnt_final_Z[3]), .FCI(tap_cnt_17_i_m2_cry_2), .S(N_77), 
        .Y(tapcnt_final_RNIES844_Y_0[3]), .FCO(tap_cnt_17_i_m2_cry_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[23]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[23]), .C(
        un10_early_flags[23]), .Y(late_flags_7_fast_0[23]));
    SLE \late_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[6])
        );
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_182  (.A(
        late_flags_Z[67]), .B(late_flags_Z[66]), .C(late_flags_Z[65]), 
        .D(late_flags_Z[64]), .Y(calc_done25_182));
    SLE \early_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[21]), 
        .D(early_flags_Z[85]), .FCI(early_flags_pmux_126_1_1_co1_5), 
        .S(early_flags_pmux_126_1_1_wmux_13_S_0), .Y(
        early_flags_pmux_126_1_1_y0_5), .FCO(
        early_flags_pmux_126_1_1_co0_6));
    SLE \tapcnt_final_upd[0]  (.D(tapcnt_final_upd_8_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[7]), .D(
        late_flags_Z[71]), .FCI(late_flags_pmux_126_1_0_co1_4), .S(
        late_flags_pmux_126_1_0_wmux_11_S_0), .Y(
        late_flags_pmux_126_1_0_y0_4), .FCO(
        late_flags_pmux_126_1_0_co0_5));
    SLE \late_flags[40]  (.D(late_flags_7_fast_0[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[40]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[30]), 
        .D(late_flags_Z[94]), .FCI(late_flags_pmux_63_1_0_co1_7), .S(
        late_flags_pmux_63_1_0_wmux_17_S_0), .Y(
        late_flags_pmux_63_1_0_y0_7), .FCO(
        late_flags_pmux_63_1_0_co0_8));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_91 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[67]), .Y(
        un10_early_flags[91]));
    SLE \early_flags[108]  (.D(early_flags_7_fast_0[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[108]));
    CFG4 #( .INIT(16'h0040) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state159  (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state155_1), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state159));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_35 (.A(
        un10_early_flags_2_0[32]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_2_Z[35]), .Y(un10_early_flags[35]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[70]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[70]), .C(
        un10_early_flags[70]), .Y(late_flags_7_fast_0[70]));
    SLE \late_flags[116]  (.D(late_flags_7_fast_0[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[116]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[9]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[9]), .C(
        un10_early_flags[9]), .Y(early_flags_7_fast_0[9]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_53 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[5]), .C(
        un10_early_flags_2_0[52]), .Y(un10_early_flags[53]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[37]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[37]), .C(
        un10_early_flags[37]), .Y(early_flags_7_fast_0[37]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_105 (.A(
        un10_early_flags_1_Z[9]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[96]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[105]));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_228  (.A(
        calc_done25_147), .B(calc_done25_146), .C(calc_done25_145), .D(
        calc_done25_144), .Y(calc_done25_228));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_6 (.A(
        early_flags_pmux_63_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[56]), .D(early_flags_Z[120]), .FCI(
        early_flags_pmux_63_1_1_co0_2), .S(
        early_flags_pmux_63_1_1_wmux_6_S_0), .Y(
        early_flags_pmux_63_1_1_y7), .FCO(
        early_flags_pmux_63_1_1_co1_2));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[5]), .D(
        late_flags_Z[69]), .FCI(late_flags_pmux_126_1_1_co1_4), .S(
        late_flags_pmux_126_1_1_wmux_11_S_0), .Y(
        late_flags_pmux_126_1_1_y0_4), .FCO(
        late_flags_pmux_126_1_1_co0_5));
    SLE \late_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[0])
        );
    CFG3 #( .INIT(8'h74) )  un1_bitalign_curr_state152 (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[0]), .C(
        bitalign_curr_state155_1), .Y(un1_bitalign_curr_state152_Z));
    SLE \tapcnt_final_upd[6]  (.D(tapcnt_final_upd_8[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[43]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[43]), .C(
        un10_early_flags[43]), .Y(late_flags_7_fast_0[43]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[17]), 
        .D(early_flags_Z[81]), .FCI(early_flags_pmux_126_1_1_co1), .S(
        early_flags_pmux_126_1_1_wmux_1_S_0), .Y(
        early_flags_pmux_126_1_1_y0_0), .FCO(
        early_flags_pmux_126_1_1_co0_0));
    CFG4 #( .INIT(16'hC505) )  \bitalign_curr_state_34_4_0_.m10  (.A(
        BIT_ALGN_OOR_0_c), .B(calc_done_Z), .C(
        bitalign_curr_state_Z[0]), .D(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(N_11));
    SLE \no_early_no_late_val_st2[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_0), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[1]));
    SLE \noearly_nolate_diff_nxt[3]  (.D(noearly_nolate_diff_nxt_8[3]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_3));
    CFG4 #( .INIT(16'h0100) )  
        \bitalign_curr_state_34_4_0_.calc_done28  (.A(un1_tapcnt_final)
        , .B(calc_done25), .C(un1_noearly_nolate_diff_start_valid), .D(
        un1_noearly_nolate_diff_nxt_valid_Z), .Y(calc_done28));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNINKIR[3]  (.A(
        late_val_Z[3]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[3]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNINKIR_0[3]));
    SLE \early_flags[6]  (.D(early_flags_7_fast_0[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[6]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_63 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[63]));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNILIIR[2]  (.A(
        late_val_Z[2]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[2]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNILIIR_0[2]));
    SLE \early_flags[75]  (.D(early_flags_7_fast_0[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[75]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_25 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_0[24]), .C(
        un10_early_flags_2_Z[21]), .Y(un10_early_flags[25]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_154  (.A(
        early_flags_Z[31]), .B(early_flags_Z[30]), .C(
        early_flags_Z[29]), .D(early_flags_Z[28]), .Y(calc_done25_154));
    SLE \early_flags[53]  (.D(early_flags_7_fast_0[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[53]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI9IJ81[4]  (.A(early_val_Z[4])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[4]), .Y(
        early_val_RNI9IJ81_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[108]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[108]), .C(
        un10_early_flags[108]), .Y(early_flags_7_fast_0[108]));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIPMIR[4]  (.A(
        late_val_Z[4]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[4]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIPMIR_0[4]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_146  (.A(
        early_flags_Z[63]), .B(early_flags_Z[62]), .C(
        early_flags_Z[61]), .D(early_flags_Z[60]), .Y(calc_done25_146));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[20]), 
        .D(early_flags_Z[84]), .FCI(early_flags_pmux_63_1_1_co1_5), .S(
        early_flags_pmux_63_1_1_wmux_13_S_0), .Y(
        early_flags_pmux_63_1_1_y0_5), .FCO(
        early_flags_pmux_63_1_1_co0_6));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[76]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[76]), .C(
        un10_early_flags[76]), .Y(early_flags_7_fast_0[76]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[101]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[101]), .C(
        un10_early_flags[101]), .Y(early_flags_7_fast_0[101]));
    CFG3 #( .INIT(8'hE4) )  \late_flags_RNO[49]  (.A(N_208), .B(
        EYE_MONITOR_LATE_net_0_0), .C(late_flags_Z[49]), .Y(
        late_flags_RNO_0[49]));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_1_wmux_20 (.A(
        early_flags_pmux_63_1_1_y0_8), .B(early_flags_pmux_63_1_1_y3_0)
        , .C(early_flags_pmux_63_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co0_9), .S(
        early_flags_pmux_63_1_1_wmux_20_S_0), .Y(
        early_flags_pmux_63_1_1_y21), .FCO(
        early_flags_pmux_63_1_1_co1_9));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_16 (.A(
        early_flags_pmux_63_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[46]), .D(early_flags_Z[110]), .FCI(
        early_flags_pmux_63_1_0_co0_7), .S(
        early_flags_pmux_63_1_0_wmux_16_S_0), .Y(
        early_flags_pmux_63_1_0_y5_0), .FCO(
        early_flags_pmux_63_1_0_co1_7));
    SLE \early_flags[109]  (.D(early_flags_7_fast_0[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[109]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_9 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_Z[8]), .C(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[9]));
    SLE \noearly_nolate_diff_start[6]  (.D(
        noearly_nolate_diff_start_7[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_6));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[22]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[22]), .C(
        un10_early_flags[22]), .Y(early_flags_7_fast_0[22]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[58]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[58]), .C(
        un10_early_flags[58]), .Y(late_flags_7_fast_0[58]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_63_1_1_co1_3), .S(
        early_flags_pmux_63_1_1_wmux_9_S_0), .Y(
        early_flags_pmux_63_1_1_wmux_9_Y_0), .FCO(
        early_flags_pmux_63_1_1_co0_4));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_90 (.A(
        un10_early_flags_1_Z[10]), .B(tap_cnt_Z[5]), .C(
        un10_early_flags_1_Z[80]), .D(un10_early_flags_2_Z[10]), .Y(
        un10_early_flags[90]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[82]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[82]), .C(
        un10_early_flags[82]), .Y(early_flags_7_fast_0[82]));
    SLE \noearly_nolate_diff_start[2]  (.D(
        noearly_nolate_diff_start_7[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_2));
    SLE \early_flags[19]  (.D(early_flags_7_fast_0[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[19]));
    SLE \late_flags[53]  (.D(late_flags_7_fast_0[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[53]));
    SLE \early_flags[20]  (.D(early_flags_7_fast_0[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[20]));
    CFG2 #( .INIT(4'hE) )  un1_bitalign_curr_state_14_1 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[1]), .Y(
        un1_bitalign_curr_state_14_1_Z));
    SLE \late_flags[90]  (.D(late_flags_7_fast_0[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[90]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[12]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[12]), .C(
        un10_early_flags[12]), .Y(late_flags_7_fast_0[12]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_171  (.A(
        late_flags_Z[35]), .B(late_flags_Z[34]), .C(late_flags_Z[33]), 
        .D(late_flags_Z[32]), .Y(calc_done25_171));
    CFG4 #( .INIT(16'hFFFE) )  
        \bitalign_curr_state_34_4_0_.un1_calc_done25_5  (.A(
        un1_tapcnt_final), .B(calc_done25), .C(
        un1_noearly_nolate_diff_start_valid), .D(
        un1_noearly_nolate_diff_nxt_valid_Z), .Y(un1_calc_done25_5));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[62]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[62]), .C(
        un10_early_flags[62]), .Y(early_flags_7_fast_0[62]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_38 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_2_0[32]), .C(
        un10_early_flags_1_Z[32]), .Y(un10_early_flags[38]));
    SLE \late_flags[85]  (.D(late_flags_7_fast_0[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[85]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[3]  (.A(VCC), .B(
        rst_cnt_Z[3]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[2]), .S(
        rst_cnt_s[3]), .Y(rst_cnt_cry_Y_1[3]), .FCO(rst_cnt_cry_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[39]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[39]), .C(
        un10_early_flags[39]), .Y(late_flags_7_fast_0[39]));
    SLE \early_flags[114]  (.D(early_flags_7_fast_0[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[114]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_1 (.A(late_val_Z[1])
        , .B(early_val_Z[1]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_0_Z), .S(tapcnt_final27_cry_1_S_0), .Y(
        tapcnt_final27_cry_1_Y_0), .FCO(tapcnt_final27_cry_1_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_7 (.A(
        early_flags_pmux_126_1_1_y7), .B(early_flags_pmux_126_1_1_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_1_co1_2), .S(
        early_flags_pmux_126_1_1_wmux_7_S_0), .Y(
        early_flags_pmux_126_1_1_y0_3), .FCO(
        early_flags_pmux_126_1_1_co0_3));
    CFG2 #( .INIT(4'h8) )  tap_cnt_0_sqmuxa_0 (.A(
        bitalign_curr_state_Z[0]), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(tap_cnt_0_sqmuxa_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[8]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[8]), .C(
        un10_early_flags[8]), .Y(late_flags_7_fast_0[8]));
    CFG4 #( .INIT(16'hA888) )  un2_early_late_diff_validlto3 (.A(
        early_late_diff_Z[3]), .B(early_late_diff_Z[2]), .C(
        early_late_diff_Z[1]), .D(early_late_diff_Z[0]), .Y(
        un2_early_late_diff_validlt7));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_5 (.A(
        un16_tapcnt_final_5), .B(un10_tapcnt_final_5), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_4_Z), .S(
        un16_tapcnt_final_cry_5_S_0), .Y(un16_tapcnt_final_cry_5_Y_0), 
        .FCO(un16_tapcnt_final_cry_5_Z));
    SLE \rst_cnt[9]  (.D(rst_cnt_s_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[9]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[29]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[29]), .C(
        un10_early_flags[29]), .Y(late_flags_7_fast_0[29]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[39]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[39]), .C(
        un10_early_flags[39]), .Y(early_flags_7_fast_0[39]));
    SLE \late_flags[15]  (.D(late_flags_7_fast_0[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[15]));
    SLE \early_flags[101]  (.D(early_flags_7_fast_0[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[101]));
    SLE \late_flags[63]  (.D(late_flags_7_fast_0[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[63]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_28 (.A(
        un10_early_flags_2_0[28]), .B(un10_early_flags_1_Z[16]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[28]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[10]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[10]), .C(
        un10_early_flags[10]), .Y(early_flags_7_fast_0[10]));
    CFG4 #( .INIT(16'hFF40) )  un1_rx_BIT_ALGN_LOAD_0_sqmuxa (.A(
        calc_done_Z), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .C(
        bitalign_curr_state154_Z), .D(rx_BIT_ALGN_LOAD_0_sqmuxa_Z), .Y(
        un1_rx_BIT_ALGN_LOAD_0_sqmuxa_i_0));
    CFG3 #( .INIT(8'h10) )  
        \bitalign_curr_state_34_4_0_.bitalign_curr_state_2_sqmuxa_4_0_0  
        (.A(bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[1]), 
        .C(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state_2_sqmuxa_4_0_0));
    CFG2 #( .INIT(4'h8) )  
        \bitalign_curr_state155.bitalign_curr_state155_1  (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state155_1));
    CFG3 #( .INIT(8'h20) )  \bitalign_curr_state_34_4_0_.m72  (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state_Z[0]), 
        .C(bitalign_curr_state61), .Y(N_116_mux));
    SLE \early_flags[22]  (.D(early_flags_7_fast_0[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[22]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[78]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[78]), .C(
        un10_early_flags[78]), .Y(late_flags_7_fast_0[78]));
    CFG2 #( .INIT(4'hE) )  un1_calc_done25_7 (.A(un1_calc_done25_5), 
        .B(un1_early_late_diff_valid_Z), .Y(un1_calc_done25_7_i));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[1]  (.A(
        tapcnt_final_13_Z[2]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[1]), .Y(tapcnt_final_13_1_Z[1]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[0]), 
        .D(early_flags_Z[64]), .FCI(VCC), .S(
        early_flags_pmux_63_1_1_wmux_S_0), .Y(
        early_flags_pmux_63_1_1_y0), .FCO(early_flags_pmux_63_1_1_co0));
    SLE \early_flags[103]  (.D(early_flags_7_fast_0[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[103]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_127 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[127]));
    SLE \late_flags[124]  (.D(late_flags_7_fast_0[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[124]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_4 (.A(late_val_Z[4])
        , .B(early_val_Z[4]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_3_Z), .S(tapcnt_final27_cry_4_S_0), .Y(
        tapcnt_final27_cry_4_Y_0), .FCO(tapcnt_final27_cry_4_Z));
    ARI1 #( .INIT(20'h45500) )  restart_trng_fg_RNIBNT7 (.A(VCC), .B(
        restart_trng_fg_i), .C(GND), .D(GND), .FCI(VCC), .S(
        restart_trng_fg_RNIBNT7_S_0), .Y(restart_trng_fg_RNIBNT7_Y_0), 
        .FCO(timeout_cnt_cry_cy));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[21]), 
        .D(late_flags_Z[85]), .FCI(late_flags_pmux_126_1_1_co1_5), .S(
        late_flags_pmux_126_1_1_wmux_13_S_0), .Y(
        late_flags_pmux_126_1_1_y0_5), .FCO(
        late_flags_pmux_126_1_1_co0_6));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[112]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[112]), .C(
        un10_early_flags[112]), .Y(late_flags_7_fast_0[112]));
    SLE \late_flags[45]  (.D(late_flags_7_fast_0[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[45]));
    CFG3 #( .INIT(8'h80) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state154_Z), 
        .C(calc_done_Z), .Y(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z));
    SLE \late_flags[28]  (.D(late_flags_7_fast_0[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[28]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_144  (.A(
        early_flags_Z[55]), .B(early_flags_Z[54]), .C(
        early_flags_Z[53]), .D(early_flags_Z[52]), .Y(calc_done25_144));
    CFG4 #( .INIT(16'h0001) )  \un1_tap_cnt_0_sqmuxa_14_i_a2[0]  (.A(
        un1_early_flags_1_sqmuxa_i), .B(N_63_0), .C(
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), .D(
        bitalign_curr_state_0_sqmuxa_10), .Y(N_89));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_3 (.A(late_val_Z[3])
        , .B(early_val_Z[3]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_2_Z), .S(tapcnt_final27_cry_3_S_0), .Y(
        tapcnt_final27_cry_3_Y_0), .FCO(tapcnt_final27_cry_3_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[36]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[36]), .C(
        un10_early_flags[36]), .Y(late_flags_7_fast_0[36]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[107]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[107]), .C(
        un10_early_flags[107]), .Y(early_flags_7_fast_0[107]));
    ARI1 #( .INIT(20'h54411) )  tapcnt_final_upd_8_cry_5_0 (.A(
        tap_cnt_Z[5]), .B(mv_dn_fg_0_sqmuxa_i_o2_0), .C(
        tapcnt_final_upd_1_sqmuxa), .D(GND), .FCI(
        tapcnt_final_upd_8_cry_4), .S(tapcnt_final_upd_8[5]), .Y(
        tapcnt_final_upd_8_cry_5_0_Y_0), .FCO(tapcnt_final_upd_8_cry_5)
        );
    CFG4 #( .INIT(16'h202F) )  \tapcnt_final_13_1_1_0[0]  (.A(
        tapcnt_final_Z[0]), .B(un1_restart_trng_fg_10_sn), .C(
        tapcnt_final_13_m0s2_0), .D(early_val_RNIBEUF3_Y[0]), .Y(
        tapcnt_final_13_1_1_0_Z[0]));
    CFG2 #( .INIT(4'h2) )  rx_BIT_ALGN_MOVE_2_sqmuxa (.A(
        un1_early_flags_1_sqmuxa_1_Z), .B(restart_trng_fg_i), .Y(
        rx_BIT_ALGN_MOVE_2_sqmuxa_Z));
    SLE \early_flags[83]  (.D(early_flags_7_fast_0[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[83]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_128  (.A(
        early_flags_Z[119]), .B(early_flags_Z[118]), .C(
        early_flags_Z[117]), .D(early_flags_Z[116]), .Y(
        calc_done25_128));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_31 (.A(
        un10_early_flags_30_0_Z), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[31]));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[5]  (.A(
        no_early_no_late_val_end1_Z[5]), .B(tapcnt_final_2_sqmuxa), .C(
        no_early_no_late_val_end2_Z[5]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[26]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[26]), .C(
        un10_early_flags[26]), .Y(late_flags_7_fast_0[26]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_s[6]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_1[0]), .C(emflag_cnt_Z[6]), .D(GND), .FCI(
        emflag_cnt_cry_Z[5]), .S(emflag_cnt_s_Z[6]), .Y(
        emflag_cnt_s_Y_0[6]), .FCO(emflag_cnt_s_FCO_0[6]));
    SLE \late_flags[118]  (.D(late_flags_7_fast_0[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[118]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_7 (.A(
        early_flags_pmux_63_1_1_y7), .B(early_flags_pmux_63_1_1_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co1_2), .S(
        early_flags_pmux_63_1_1_wmux_7_S_0), .Y(
        early_flags_pmux_63_1_1_y0_3), .FCO(
        early_flags_pmux_63_1_1_co0_3));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[28]), 
        .D(early_flags_Z[92]), .FCI(early_flags_pmux_63_1_1_co1_7), .S(
        early_flags_pmux_63_1_1_wmux_17_S_0), .Y(
        early_flags_pmux_63_1_1_y0_7), .FCO(
        early_flags_pmux_63_1_1_co0_8));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[126]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[126]), .C(
        un10_early_flags[126]), .Y(early_flags_7_fast_0[126]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_6_0 (.A(
        emflag_cnt_Z[6]), .B(un1_restart_trng_fg_5_0), .C(
        no_early_no_late_val_st2_Z[6]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_5), .S(
        noearly_nolate_diff_nxt_8[6]), .Y(
        noearly_nolate_diff_nxt_8_cry_6_0_Y_0), .FCO(
        noearly_nolate_diff_nxt_8_cry_6));
    CFG4 #( .INIT(16'h8000) )  
        \bitalign_curr_state_34_4_0_.calc_done25_227  (.A(
        calc_done25_143), .B(calc_done25_142), .C(calc_done25_141), .D(
        calc_done25_140), .Y(calc_done25_227));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_4 (.A(
        early_flags_pmux_126_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[41]), .D(early_flags_Z[105]), .FCI(
        early_flags_pmux_126_1_1_co0_1), .S(
        early_flags_pmux_126_1_1_wmux_4_S_0), .Y(
        early_flags_pmux_126_1_1_y5), .FCO(
        early_flags_pmux_126_1_1_co1_1));
    CFG3 #( .INIT(8'h40) )  rx_trng_done_RNO (.A(restart_trng_fg_i), 
        .B(bitalign_curr_state41_Z), .C(bitalign_curr_state_Z[1]), .Y(
        N_1403));
    CFG4 #( .INIT(16'hF1F0) )  rx_trng_done_0_sqmuxa_i (.A(
        early_flags_1_sqmuxa_1_Z), .B(un1_bitalign_curr_state_13_1_Z), 
        .C(restart_trng_fg_i), .D(un1_bitalign_curr_state148_2_Z), .Y(
        rx_trng_done_0_sqmuxa_i_Z));
    SLE \late_flags[78]  (.D(late_flags_7_fast_0[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[78]));
    SLE \no_early_no_late_val_end1[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[3]));
    CFG4 #( .INIT(16'h0001) )  
        \bitalign_curr_state_34_4_0_.calc_done25_173  (.A(
        late_flags_Z[59]), .B(late_flags_Z[58]), .C(late_flags_Z[57]), 
        .D(late_flags_Z[56]), .Y(calc_done25_173));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_30_0 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[6]), .Y(un10_early_flags_30_0_Z));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIJ5QFH[4]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIPMIR_0[4]), .B(
        early_val_RNI9IJ81_Z[4]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[4]), .FCI(tapcnt_final_13_m1_cry_3), .S(
        tapcnt_final_13_m1[4]), .Y(early_val_RNIJ5QFH_Y[4]), .FCO(
        tapcnt_final_13_m1_cry_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[14]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[14]), .C(
        un10_early_flags[14]), .Y(early_flags_7_fast_0[14]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_21 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[16]), .C(
        un10_early_flags_2_Z[21]), .Y(un10_early_flags[21]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[18]), 
        .D(late_flags_Z[82]), .FCI(late_flags_pmux_63_1_0_0_co1), .S(
        late_flags_pmux_63_1_0_wmux_1_S_0), .Y(
        late_flags_pmux_63_1_0_y0_0), .FCO(
        late_flags_pmux_63_1_0_co0_0));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_127_1_0_wmux (.A(
        emflag_cnt_Z[1]), .B(emflag_cnt_Z[0]), .C(
        early_flags_pmux_63_1_1_wmux_10_Y_0), .D(
        early_flags_pmux_63_1_0_wmux_10_Y_0), .FCI(VCC), .S(
        early_flags_pmux_127_1_0_wmux_S_0), .Y(
        early_flags_pmux_127_1_0_y0), .FCO(
        early_flags_pmux_127_1_0_co0));
    
endmodule


module 
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_0s_0s_0s_26s_10s_10s_0(
        
       EYE_MONITOR_LATE_net_0_0,
       EYE_MONITOR_EARLY_net_0_0,
       BIT_ALGN_EYE_IN_c,
       RX_CLK_ALIGN_DONE_arst,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       debouncer_0_DB_OUT,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE,
       BIT_ALGN_ERR_c,
       BIT_ALGN_OOR_0_c,
       BIT_ALGN_START_0_c,
       BIT_ALGN_DONE_0_c,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS,
       PLL_LOCK_0
    );
input  EYE_MONITOR_LATE_net_0_0;
input  EYE_MONITOR_EARLY_net_0_0;
input  [2:0] BIT_ALGN_EYE_IN_c;
input  RX_CLK_ALIGN_DONE_arst;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  debouncer_0_DB_OUT;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE;
output BIT_ALGN_ERR_c;
input  BIT_ALGN_OOR_0_c;
output BIT_ALGN_START_0_c;
output BIT_ALGN_DONE_0_c;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS;
input  PLL_LOCK_0;

    wire GND, VCC;
    
    
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_TRNG_Z1_0 
        u_CoreRxIODBitAlign (.BIT_ALGN_EYE_IN_c({BIT_ALGN_EYE_IN_c[2], 
        BIT_ALGN_EYE_IN_c[1], BIT_ALGN_EYE_IN_c[0]}), 
        .EYE_MONITOR_EARLY_net_0_0(EYE_MONITOR_EARLY_net_0_0), 
        .EYE_MONITOR_LATE_net_0_0(EYE_MONITOR_LATE_net_0_0), 
        .PLL_LOCK_0(PLL_LOCK_0), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS), .BIT_ALGN_DONE_0_c(
        BIT_ALGN_DONE_0_c), .BIT_ALGN_START_0_c(BIT_ALGN_START_0_c), 
        .BIT_ALGN_OOR_0_c(BIT_ALGN_OOR_0_c), .BIT_ALGN_ERR_c(
        BIT_ALGN_ERR_c), .CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module CORERXIODBITALIGN_C0_1(
       BIT_ALGN_EYE_IN_c,
       EYE_MONITOR_EARLY_net_0_0,
       EYE_MONITOR_LATE_net_0_0,
       PLL_LOCK_0,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS,
       BIT_ALGN_DONE_0_c,
       BIT_ALGN_START_0_c,
       BIT_ALGN_OOR_0_c,
       BIT_ALGN_ERR_c,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD,
       debouncer_0_DB_OUT,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst
    );
input  [2:0] BIT_ALGN_EYE_IN_c;
input  EYE_MONITOR_EARLY_net_0_0;
input  EYE_MONITOR_LATE_net_0_0;
input  PLL_LOCK_0;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS;
output BIT_ALGN_DONE_0_c;
output BIT_ALGN_START_0_c;
input  BIT_ALGN_OOR_0_c;
output BIT_ALGN_ERR_c;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR;
output CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD;
input  debouncer_0_DB_OUT;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  RX_CLK_ALIGN_DONE_arst;

    wire GND, VCC;
    
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_0s_0s_0s_26s_10s_10s_0 
        CORERXIODBITALIGN_C0_0 (.EYE_MONITOR_LATE_net_0_0(
        EYE_MONITOR_LATE_net_0_0), .EYE_MONITOR_EARLY_net_0_0(
        EYE_MONITOR_EARLY_net_0_0), .BIT_ALGN_EYE_IN_c({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE), .BIT_ALGN_ERR_c(
        BIT_ALGN_ERR_c), .BIT_ALGN_OOR_0_c(BIT_ALGN_OOR_0_c), 
        .BIT_ALGN_START_0_c(BIT_ALGN_START_0_c), .BIT_ALGN_DONE_0_c(
        BIT_ALGN_DONE_0_c), .CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS), .PLL_LOCK_0(
        PLL_LOCK_0));
    
endmodule


module PF_OSC_C1_PF_OSC_C1_0_PF_OSC(
       PF_OSC_C1_0_RCOSC_160MHZ_GL
    );
output PF_OSC_C1_0_RCOSC_160MHZ_GL;

    wire I_OSC_160_CLK_c, VCC, GND;
    
    VCC VCC_Z (.Y(VCC));
    OSC_RC160MHZ I_OSC_160 (.OSC_160MHZ_ON(VCC), .CLK(I_OSC_160_CLK_c));
    CLKINT I_OSC_160_INT (.A(I_OSC_160_CLK_c), .Y(
        PF_OSC_C1_0_RCOSC_160MHZ_GL));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_OSC_C1(
       PF_OSC_C1_0_RCOSC_160MHZ_GL
    );
output PF_OSC_C1_0_RCOSC_160MHZ_GL;

    wire GND, VCC;
    
    PF_OSC_C1_PF_OSC_C1_0_PF_OSC PF_OSC_C1_0 (
        .PF_OSC_C1_0_RCOSC_160MHZ_GL(PF_OSC_C1_0_RCOSC_160MHZ_GL));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_TX_C0_PF_IOD_TX_CLK_PF_IOD(
       TX_CLK,
       TX_CLK_N,
       LANECTRL_ADDR_CMD_0_TX_DQS_270,
       LANECTRL_ADDR_CMD_0_TX_DQS,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90,
       LANECTRL_ADDR_CMD_0_TX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_RX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_ARST_N,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G
    );
output TX_CLK;
output TX_CLK_N;
input  LANECTRL_ADDR_CMD_0_TX_DQS_270;
input  LANECTRL_ADDR_CMD_0_TX_DQS;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90;
input  LANECTRL_ADDR_CMD_0_TX_SYNC_RST;
input  LANECTRL_ADDR_CMD_0_RX_SYNC_RST;
input  LANECTRL_ADDR_CMD_0_ARST_N;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;

    wire [1:0] RX_DATA_4;
    wire [9:2] RX_DATA_2;
    wire [10:0] CDR_CLK_B_SEL_4;
    wire VCC, GND, EYE_MONITOR_EARLY_1, EYE_MONITOR_LATE_1, 
        DELAY_LINE_OUT_OF_RANGE_5, D_I_OUTBUF_DIFF_0_net, OE_4, 
        DDR_DO_READ_4, CDR_CLK_A_SEL_8_4, CDR_CLK_A_SEL_9_4, 
        CDR_CLK_A_SEL_10_4, SWITCH_5, CDR_CLR_NEXT_CLK_N_4, 
        TX_DATA_OUT_9_4, TX_DATA_OUT_8_4, AL_N_OUT_4, OUTFF_SL_OUT_4, 
        OUTFF_EN_OUT_4, INFF_SL_OUT_4, INFF_EN_OUT_4, RX_CLK_OUT_4, 
        TX_CLK_OUT_4;
    
    OUTBUF_DIFF I_OUTBUF_DIFF_0 (.D(D_I_OUTBUF_DIFF_0_net), .PADP(
        TX_CLK), .PADN(TX_CLK_N));
    VCC VCC_Z (.Y(VCC));
    IOD #( .DATA_RATE(1000.000000), .FORMAL_NAME("TX_CLK"), .INTERFACE_NAME("TX_DDRX_B_C")
        , .DELAY_LINE_SIMULATION_MODE("DISABLED"), .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000)
        , .RESERVED_0(1'b0), .RX_CLK_EN(1'b0), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b1)
        , .TX_CLK_INV(1'b0), .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b10), .RX_MODE(4'b0000), .EYE_MONITOR_MODE(1'b0)
        , .DYN_DELAY_LINE_EN(1'b0), .FIFO_WR_EN(1'b0), .EYE_MONITOR_EN(1'b0)
        , .TX_MODE(7'b1000010), .TX_CLK_SEL(2'b10), .TX_OE_MODE(3'b010)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b0)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b0)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b00)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_0 (.EYE_MONITOR_EARLY(EYE_MONITOR_EARLY_1), 
        .EYE_MONITOR_LATE(EYE_MONITOR_LATE_1), .RX_DATA({RX_DATA_2[9], 
        RX_DATA_2[8], RX_DATA_2[7], RX_DATA_2[6], RX_DATA_2[5], 
        RX_DATA_2[4], RX_DATA_2[3], RX_DATA_2[2], RX_DATA_4[1], 
        RX_DATA_4[0]}), .DELAY_LINE_OUT_OF_RANGE(
        DELAY_LINE_OUT_OF_RANGE_5), .TX_DATA({GND, GND, GND, GND, GND, 
        VCC, GND, VCC}), .OE_DATA({GND, GND, VCC, VCC}), .RX_BIT_SLIP(
        GND), .EYE_MONITOR_CLEAR_FLAGS(GND), .DELAY_LINE_MOVE(GND), 
        .DELAY_LINE_DIRECTION(GND), .DELAY_LINE_LOAD(GND), .RX_CLK(GND)
        , .TX_CLK(PF_IOD_TX_CCC_C0_0_TX_CLK_G), .ODT_EN(GND), .INFF_SL(
        GND), .INFF_EN(GND), .OUTFF_SL(GND), .OUTFF_EN(GND), .AL_N(GND)
        , .OEFF_LAT_N(GND), .OEFF_SD_N(GND), .OEFF_AD_N(GND), 
        .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(GND), 
        .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), .RX_P(
        GND), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(GND), .ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, 
        GND, GND, PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90}), 
        .RX_DQS_90({GND, GND}), .TX_DQS(LANECTRL_ADDR_CMD_0_TX_DQS), 
        .TX_DQS_270(LANECTRL_ADDR_CMD_0_TX_DQS_270), .FIFO_WR_PTR({GND, 
        GND, GND}), .FIFO_RD_PTR({GND, GND, GND}), .TX(
        D_I_OUTBUF_DIFF_0_net), .OE(OE_4), .CDR_CLK(GND), 
        .CDR_NEXT_CLK(GND), .EYE_MONITOR_LANE_WIDTH({GND, GND, GND}), 
        .DDR_DO_READ(DDR_DO_READ_4), .CDR_CLK_A_SEL_8(
        CDR_CLK_A_SEL_8_4), .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9_4), 
        .CDR_CLK_A_SEL_10(CDR_CLK_A_SEL_10_4), .CDR_CLK_B_SEL({
        CDR_CLK_B_SEL_4[10], CDR_CLK_B_SEL_4[9], CDR_CLK_B_SEL_4[8], 
        CDR_CLK_B_SEL_4[7], CDR_CLK_B_SEL_4[6], CDR_CLK_B_SEL_4[5], 
        CDR_CLK_B_SEL_4[4], CDR_CLK_B_SEL_4[3], CDR_CLK_B_SEL_4[2], 
        CDR_CLK_B_SEL_4[1], CDR_CLK_B_SEL_4[0]}), .SWITCH(SWITCH_5), 
        .CDR_CLR_NEXT_CLK_N(CDR_CLR_NEXT_CLK_N_4), .TX_DATA_OUT_9(
        TX_DATA_OUT_9_4), .TX_DATA_OUT_8(TX_DATA_OUT_8_4), .AL_N_OUT(
        AL_N_OUT_4), .OUTFF_SL_OUT(OUTFF_SL_OUT_4), .OUTFF_EN_OUT(
        OUTFF_EN_OUT_4), .INFF_SL_OUT(INFF_SL_OUT_4), .INFF_EN_OUT(
        INFF_EN_OUT_4), .RX_CLK_OUT(RX_CLK_OUT_4), .TX_CLK_OUT(
        TX_CLK_OUT_4));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_TX_C0_PF_IOD_TX_PF_IOD(
       TXD,
       TXD_N,
       prbsgen_parallel_fab_0_prbs_out_msb_o_0,
       LANECTRL_ADDR_CMD_0_TX_DQS_270,
       LANECTRL_ADDR_CMD_0_TX_DQS,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0,
       LANECTRL_ADDR_CMD_0_TX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_RX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_ARST_N,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G
    );
output [1:0] TXD;
output [1:0] TXD_N;
input  [7:0] prbsgen_parallel_fab_0_prbs_out_msb_o_0;
input  LANECTRL_ADDR_CMD_0_TX_DQS_270;
input  LANECTRL_ADDR_CMD_0_TX_DQS;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0;
input  LANECTRL_ADDR_CMD_0_TX_SYNC_RST;
input  LANECTRL_ADDR_CMD_0_RX_SYNC_RST;
input  LANECTRL_ADDR_CMD_0_ARST_N;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;

    wire [1:0] RX_DATA_2;
    wire [9:2] RX_DATA_0;
    wire [10:0] CDR_CLK_B_SEL_2;
    wire [1:0] RX_DATA_3;
    wire [9:2] RX_DATA_1;
    wire [10:0] CDR_CLK_B_SEL_3;
    wire VCC, GND, EYE_MONITOR_EARLY, EYE_MONITOR_LATE, 
        DELAY_LINE_OUT_OF_RANGE_3, D_I_OUTBUF_DIFF_0_net, OE_2, 
        DDR_DO_READ_2, CDR_CLK_A_SEL_8_2, CDR_CLK_A_SEL_9_2, 
        CDR_CLK_A_SEL_10_2, SWITCH_3, CDR_CLR_NEXT_CLK_N_2, 
        TX_DATA_OUT_9_2, TX_DATA_OUT_8_2, AL_N_OUT_2, OUTFF_SL_OUT_2, 
        OUTFF_EN_OUT_2, INFF_SL_OUT_2, INFF_EN_OUT_2, RX_CLK_OUT_2, 
        TX_CLK_OUT_2, D_I_OUTBUF_DIFF_1_net, EYE_MONITOR_EARLY_0, 
        EYE_MONITOR_LATE_0, DELAY_LINE_OUT_OF_RANGE_4, OE_3, 
        DDR_DO_READ_3, CDR_CLK_A_SEL_8_3, CDR_CLK_A_SEL_9_3, 
        CDR_CLK_A_SEL_10_3, SWITCH_4, CDR_CLR_NEXT_CLK_N_3, 
        TX_DATA_OUT_9_3, TX_DATA_OUT_8_3, AL_N_OUT_3, OUTFF_SL_OUT_3, 
        OUTFF_EN_OUT_3, INFF_SL_OUT_3, INFF_EN_OUT_3, RX_CLK_OUT_3, 
        TX_CLK_OUT_3;
    
    OUTBUF_DIFF I_OUTBUF_DIFF_0 (.D(D_I_OUTBUF_DIFF_0_net), .PADP(
        TXD[0]), .PADN(TXD_N[0]));
    IOD #( .DATA_RATE(1000.000000), .FORMAL_NAME("TXD"), .INTERFACE_NAME("TX_DDRX_B_C")
        , .DELAY_LINE_SIMULATION_MODE("DISABLED"), .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000)
        , .RESERVED_0(1'b0), .RX_CLK_EN(1'b0), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b1)
        , .TX_CLK_INV(1'b0), .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b10), .RX_MODE(4'b0000), .EYE_MONITOR_MODE(1'b0)
        , .DYN_DELAY_LINE_EN(1'b0), .FIFO_WR_EN(1'b0), .EYE_MONITOR_EN(1'b0)
        , .TX_MODE(7'b1000100), .TX_CLK_SEL(2'b11), .TX_OE_MODE(3'b010)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b0)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b0)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b00)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_1 (.EYE_MONITOR_EARLY(EYE_MONITOR_EARLY_0), 
        .EYE_MONITOR_LATE(EYE_MONITOR_LATE_0), .RX_DATA({RX_DATA_1[9], 
        RX_DATA_1[8], RX_DATA_1[7], RX_DATA_1[6], RX_DATA_1[5], 
        RX_DATA_1[4], RX_DATA_1[3], RX_DATA_1[2], RX_DATA_3[1], 
        RX_DATA_3[0]}), .DELAY_LINE_OUT_OF_RANGE(
        DELAY_LINE_OUT_OF_RANGE_4), .TX_DATA({
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[0]}), .OE_DATA({VCC, 
        VCC, VCC, VCC}), .RX_BIT_SLIP(GND), .EYE_MONITOR_CLEAR_FLAGS(
        GND), .DELAY_LINE_MOVE(GND), .DELAY_LINE_DIRECTION(GND), 
        .DELAY_LINE_LOAD(GND), .RX_CLK(GND), .TX_CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .ODT_EN(GND), .INFF_SL(GND), 
        .INFF_EN(GND), .OUTFF_SL(GND), .OUTFF_EN(GND), .AL_N(GND), 
        .OEFF_LAT_N(GND), .OEFF_SD_N(GND), .OEFF_AD_N(GND), 
        .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(GND), 
        .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), .RX_P(
        GND), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(GND), .ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, 
        GND, GND, PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0}), 
        .RX_DQS_90({GND, GND}), .TX_DQS(LANECTRL_ADDR_CMD_0_TX_DQS), 
        .TX_DQS_270(LANECTRL_ADDR_CMD_0_TX_DQS_270), .FIFO_WR_PTR({GND, 
        GND, GND}), .FIFO_RD_PTR({GND, GND, GND}), .TX(
        D_I_OUTBUF_DIFF_1_net), .OE(OE_3), .CDR_CLK(GND), 
        .CDR_NEXT_CLK(GND), .EYE_MONITOR_LANE_WIDTH({GND, GND, GND}), 
        .DDR_DO_READ(DDR_DO_READ_3), .CDR_CLK_A_SEL_8(
        CDR_CLK_A_SEL_8_3), .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9_3), 
        .CDR_CLK_A_SEL_10(CDR_CLK_A_SEL_10_3), .CDR_CLK_B_SEL({
        CDR_CLK_B_SEL_3[10], CDR_CLK_B_SEL_3[9], CDR_CLK_B_SEL_3[8], 
        CDR_CLK_B_SEL_3[7], CDR_CLK_B_SEL_3[6], CDR_CLK_B_SEL_3[5], 
        CDR_CLK_B_SEL_3[4], CDR_CLK_B_SEL_3[3], CDR_CLK_B_SEL_3[2], 
        CDR_CLK_B_SEL_3[1], CDR_CLK_B_SEL_3[0]}), .SWITCH(SWITCH_4), 
        .CDR_CLR_NEXT_CLK_N(CDR_CLR_NEXT_CLK_N_3), .TX_DATA_OUT_9(
        TX_DATA_OUT_9_3), .TX_DATA_OUT_8(TX_DATA_OUT_8_3), .AL_N_OUT(
        AL_N_OUT_3), .OUTFF_SL_OUT(OUTFF_SL_OUT_3), .OUTFF_EN_OUT(
        OUTFF_EN_OUT_3), .INFF_SL_OUT(INFF_SL_OUT_3), .INFF_EN_OUT(
        INFF_EN_OUT_3), .RX_CLK_OUT(RX_CLK_OUT_3), .TX_CLK_OUT(
        TX_CLK_OUT_3));
    VCC VCC_Z (.Y(VCC));
    OUTBUF_DIFF I_OUTBUF_DIFF_1 (.D(D_I_OUTBUF_DIFF_1_net), .PADP(
        TXD[1]), .PADN(TXD_N[1]));
    IOD #( .DATA_RATE(1000.000000), .FORMAL_NAME("TXD:NO_IOD_N_SIDE")
        , .INTERFACE_NAME("TX_DDRX_B_C"), .DELAY_LINE_SIMULATION_MODE("DISABLED")
        , .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000), .RESERVED_0(1'b0)
        , .RX_CLK_EN(1'b0), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b1), .TX_CLK_INV(1'b0)
        , .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b10), .RX_MODE(4'b0000), .EYE_MONITOR_MODE(1'b0)
        , .DYN_DELAY_LINE_EN(1'b0), .FIFO_WR_EN(1'b0), .EYE_MONITOR_EN(1'b0)
        , .TX_MODE(7'b1000100), .TX_CLK_SEL(2'b11), .TX_OE_MODE(3'b010)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b0)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b0)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b00)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_0 (.EYE_MONITOR_EARLY(EYE_MONITOR_EARLY), 
        .EYE_MONITOR_LATE(EYE_MONITOR_LATE), .RX_DATA({RX_DATA_0[9], 
        RX_DATA_0[8], RX_DATA_0[7], RX_DATA_0[6], RX_DATA_0[5], 
        RX_DATA_0[4], RX_DATA_0[3], RX_DATA_0[2], RX_DATA_2[1], 
        RX_DATA_2[0]}), .DELAY_LINE_OUT_OF_RANGE(
        DELAY_LINE_OUT_OF_RANGE_3), .TX_DATA({
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[0]}), .OE_DATA({VCC, 
        VCC, VCC, VCC}), .RX_BIT_SLIP(GND), .EYE_MONITOR_CLEAR_FLAGS(
        GND), .DELAY_LINE_MOVE(GND), .DELAY_LINE_DIRECTION(GND), 
        .DELAY_LINE_LOAD(GND), .RX_CLK(GND), .TX_CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .ODT_EN(GND), .INFF_SL(GND), 
        .INFF_EN(GND), .OUTFF_SL(GND), .OUTFF_EN(GND), .AL_N(GND), 
        .OEFF_LAT_N(GND), .OEFF_SD_N(GND), .OEFF_AD_N(GND), 
        .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(GND), 
        .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), .RX_P(
        GND), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(GND), .ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, 
        GND, GND, PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0}), 
        .RX_DQS_90({GND, GND}), .TX_DQS(LANECTRL_ADDR_CMD_0_TX_DQS), 
        .TX_DQS_270(LANECTRL_ADDR_CMD_0_TX_DQS_270), .FIFO_WR_PTR({GND, 
        GND, GND}), .FIFO_RD_PTR({GND, GND, GND}), .TX(
        D_I_OUTBUF_DIFF_0_net), .OE(OE_2), .CDR_CLK(GND), 
        .CDR_NEXT_CLK(GND), .EYE_MONITOR_LANE_WIDTH({GND, GND, GND}), 
        .DDR_DO_READ(DDR_DO_READ_2), .CDR_CLK_A_SEL_8(
        CDR_CLK_A_SEL_8_2), .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9_2), 
        .CDR_CLK_A_SEL_10(CDR_CLK_A_SEL_10_2), .CDR_CLK_B_SEL({
        CDR_CLK_B_SEL_2[10], CDR_CLK_B_SEL_2[9], CDR_CLK_B_SEL_2[8], 
        CDR_CLK_B_SEL_2[7], CDR_CLK_B_SEL_2[6], CDR_CLK_B_SEL_2[5], 
        CDR_CLK_B_SEL_2[4], CDR_CLK_B_SEL_2[3], CDR_CLK_B_SEL_2[2], 
        CDR_CLK_B_SEL_2[1], CDR_CLK_B_SEL_2[0]}), .SWITCH(SWITCH_3), 
        .CDR_CLR_NEXT_CLK_N(CDR_CLR_NEXT_CLK_N_2), .TX_DATA_OUT_9(
        TX_DATA_OUT_9_2), .TX_DATA_OUT_8(TX_DATA_OUT_8_2), .AL_N_OUT(
        AL_N_OUT_2), .OUTFF_SL_OUT(OUTFF_SL_OUT_2), .OUTFF_EN_OUT(
        OUTFF_EN_OUT_2), .INFF_SL_OUT(INFF_SL_OUT_2), .INFF_EN_OUT(
        INFF_EN_OUT_2), .RX_CLK_OUT(RX_CLK_OUT_2), .TX_CLK_OUT(
        TX_CLK_OUT_2));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_TX_C0_PF_IOD_CLK_TRAINING_PF_IOD(
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0,
       LANECTRL_ADDR_CMD_0_TX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_RX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_ARST_N,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G
    );
output [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0;
input  LANECTRL_ADDR_CMD_0_TX_SYNC_RST;
input  LANECTRL_ADDR_CMD_0_RX_SYNC_RST;
input  LANECTRL_ADDR_CMD_0_ARST_N;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;

    wire [1:0] RX_DATA_5;
    wire [7:1] RX_DATA_0_net_0;
    wire [10:0] CDR_CLK_B_SEL_5;
    wire GND, VCC, EYE_MONITOR_EARLY_2, EYE_MONITOR_LATE_2, 
        DELAY_LINE_OUT_OF_RANGE_6, TX_2, OE_5, DDR_DO_READ_5, 
        CDR_CLK_A_SEL_8_5, CDR_CLK_A_SEL_9_5, CDR_CLK_A_SEL_10_5, 
        SWITCH_6, CDR_CLR_NEXT_CLK_N_5, TX_DATA_OUT_9_5, 
        TX_DATA_OUT_8_5, AL_N_OUT_5, OUTFF_SL_OUT_5, OUTFF_EN_OUT_5, 
        INFF_SL_OUT_5, INFF_EN_OUT_5, RX_CLK_OUT_5, TX_CLK_OUT_5;
    
    VCC VCC_Z (.Y(VCC));
    IOD #( .DATA_RATE(1000.000000), .FORMAL_NAME("HS_IO_CLK_TRAINING")
        , .INTERFACE_NAME("TX_DDRX_B_C"), .DELAY_LINE_SIMULATION_MODE("DISABLED")
        , .MSC_UNIQUE(""), .INTERFACE_LEVEL(3'b000), .RESERVED_0(1'b0)
        , .RX_CLK_EN(1'b1), .RX_CLK_INV(1'b0), .TX_CLK_EN(1'b0), .TX_CLK_INV(1'b0)
        , .HS_IO_CLK_SEL(3'b000), .QDR_EN(1'b0), .EDGE_DETECT_EN(1'b0)
        , .DELAY_LINE_MODE(2'b00), .RX_MODE(4'b0100), .EYE_MONITOR_MODE(1'b1)
        , .DYN_DELAY_LINE_EN(1'b0), .FIFO_WR_EN(1'b0), .EYE_MONITOR_EN(1'b1)
        , .TX_MODE(7'b0000000), .TX_CLK_SEL(2'b00), .TX_OE_MODE(3'b111)
        , .TX_OE_CLK_INV(1'b0), .RX_DELAY_VAL(7'b0000001), .RX_DELAY_VAL_X2(1'b0)
        , .TX_DELAY_VAL(7'b0000001), .EYE_MONITOR_WIDTH(3'b001), .EYE_MONITOR_WIDTH_SRC(1'b1)
        , .RESERVED_1(1'b0), .DISABLE_LANECTRL_RESET(1'b0), .INPUT_DELAY_SEL(2'b11)
        , .OEFF_EN_INV(1'b0), .INFF_EN_INV(1'b0), .OUTFF_EN_INV(1'b0)
         )  I_IOD_0 (.EYE_MONITOR_EARLY(EYE_MONITOR_EARLY_2), 
        .EYE_MONITOR_LATE(EYE_MONITOR_LATE_2), .RX_DATA({
        RX_DATA_0_net_0[7], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        RX_DATA_0_net_0[5], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        RX_DATA_0_net_0[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        RX_DATA_0_net_0[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0], 
        RX_DATA_5[1], RX_DATA_5[0]}), .DELAY_LINE_OUT_OF_RANGE(
        DELAY_LINE_OUT_OF_RANGE_6), .TX_DATA({GND, GND, GND, GND, GND, 
        GND, GND, GND}), .OE_DATA({GND, GND, GND, GND}), .RX_BIT_SLIP(
        GND), .EYE_MONITOR_CLEAR_FLAGS(VCC), .DELAY_LINE_MOVE(GND), 
        .DELAY_LINE_DIRECTION(GND), .DELAY_LINE_LOAD(GND), .RX_CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .TX_CLK(GND), .ODT_EN(GND), 
        .INFF_SL(GND), .INFF_EN(GND), .OUTFF_SL(GND), .OUTFF_EN(GND), 
        .AL_N(GND), .OEFF_LAT_N(GND), .OEFF_SD_N(GND), .OEFF_AD_N(GND), 
        .INFF_LAT_N(GND), .INFF_SD_N(GND), .INFF_AD_N(GND), 
        .OUTFF_LAT_N(GND), .OUTFF_SD_N(GND), .OUTFF_AD_N(GND), .RX_P(
        GND), .RX_N(GND), .TX_DATA_9(GND), .TX_DATA_8(GND), .ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), .HS_IO_CLK({GND, GND, GND, 
        GND, GND, PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0}), 
        .RX_DQS_90({GND, GND}), .TX_DQS(GND), .TX_DQS_270(GND), 
        .FIFO_WR_PTR({GND, GND, GND}), .FIFO_RD_PTR({GND, GND, GND}), 
        .TX(TX_2), .OE(OE_5), .CDR_CLK(GND), .CDR_NEXT_CLK(GND), 
        .EYE_MONITOR_LANE_WIDTH({GND, GND, GND}), .DDR_DO_READ(
        DDR_DO_READ_5), .CDR_CLK_A_SEL_8(CDR_CLK_A_SEL_8_5), 
        .CDR_CLK_A_SEL_9(CDR_CLK_A_SEL_9_5), .CDR_CLK_A_SEL_10(
        CDR_CLK_A_SEL_10_5), .CDR_CLK_B_SEL({CDR_CLK_B_SEL_5[10], 
        CDR_CLK_B_SEL_5[9], CDR_CLK_B_SEL_5[8], CDR_CLK_B_SEL_5[7], 
        CDR_CLK_B_SEL_5[6], CDR_CLK_B_SEL_5[5], CDR_CLK_B_SEL_5[4], 
        CDR_CLK_B_SEL_5[3], CDR_CLK_B_SEL_5[2], CDR_CLK_B_SEL_5[1], 
        CDR_CLK_B_SEL_5[0]}), .SWITCH(SWITCH_6), .CDR_CLR_NEXT_CLK_N(
        CDR_CLR_NEXT_CLK_N_5), .TX_DATA_OUT_9(TX_DATA_OUT_9_5), 
        .TX_DATA_OUT_8(TX_DATA_OUT_8_5), .AL_N_OUT(AL_N_OUT_5), 
        .OUTFF_SL_OUT(OUTFF_SL_OUT_5), .OUTFF_EN_OUT(OUTFF_EN_OUT_5), 
        .INFF_SL_OUT(INFF_SL_OUT_5), .INFF_EN_OUT(INFF_EN_OUT_5), 
        .RX_CLK_OUT(RX_CLK_OUT_5), .TX_CLK_OUT(TX_CLK_OUT_5));
    GND GND_Z (.Y(GND));
    
endmodule


module 
        PF_IOD_GENERIC_TX_C0_LANECTRL_ADDR_CMD_0_PF_LANECTRL_PAUSE_SYNC_1(
        
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net,
       OR2_PAUSE_Y
    );
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;
output HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net;
input  OR2_PAUSE_Y;

    wire VCC, pause_sync_0_i, GND;
    
    SLE \pipe.pause_sync  (.D(pause_sync_0_i), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(VCC), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net));
    VCC VCC_Z (.Y(VCC));
    SLE \pipe.pause_sync_0  (.D(OR2_PAUSE_Y), .CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .EN(VCC), .ALn(VCC), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(pause_sync_0_i));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_TX_C0_LANECTRL_ADDR_CMD_0_PF_LANECTRL(
       OR2_PAUSE_Y,
       LANECTRL_ADDR_CMD_0_TX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_RX_SYNC_RST,
       LANECTRL_ADDR_CMD_0_ARST_N,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       LANECTRL_ADDR_CMD_0_TX_DQS_270,
       LANECTRL_ADDR_CMD_0_TX_DQS
    );
input  OR2_PAUSE_Y;
output LANECTRL_ADDR_CMD_0_TX_SYNC_RST;
output LANECTRL_ADDR_CMD_0_RX_SYNC_RST;
output LANECTRL_ADDR_CMD_0_ARST_N;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;
output LANECTRL_ADDR_CMD_0_TX_DQS_270;
output LANECTRL_ADDR_CMD_0_TX_DQS;

    wire [2:0] EYE_MONITOR_WIDTH_OUT;
    wire [0:0] RX_DQS_90;
    wire [1:1] RX_DQS_90_0;
    wire [2:0] FIFO_WR_PTR;
    wire [2:0] FIFO_RD_PTR;
    wire TX_DQS, TX_DQS_270, GND, VCC, 
        HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net, RX_DATA_VALID, 
        RX_BURST_DETECT, RX_DELAY_LINE_OUT_OF_RANGE, 
        TX_DELAY_LINE_OUT_OF_RANGE, CLK_OUT_R_0, A_OUT_RST_N, 
        ODT_EN_SEL_0, CDR_CLK_0, CDR_NEXT_CLK_0, ODT_EN_OUT_0;
    
    LANECTRL #( .DATA_RATE(1000.000000), .FORMAL_NAME("LANE_RESET%DUPLICATE")
        , .INTERFACE_NAME("TX_DDRX_B_C"), .DELAY_LINE_SIMULATION_MODE("DISABLED")
        , .INTERFACE_LEVEL(3'b000), .RESERVED_0(1'b0), .RESERVED_1(1'b0)
        , .RESERVED_2(1'b0), .SOFTRESET_EN(1'b0), .SOFTRESET(1'b0), .RX_DQS_DELAY_LINE_EN(1'b0)
        , .TX_DQS_DELAY_LINE_EN(1'b1), .RX_DQS_DELAY_LINE_DIRECTION(1'b1)
        , .TX_DQS_DELAY_LINE_DIRECTION(1'b1), .RX_DQS_DELAY_VAL(8'b00000001)
        , .TX_DQS_DELAY_VAL(8'b00000001), .FIFO_EN(1'b1), .FIFO_MODE(1'b0)
        , .FIFO_RD_PTR_MODE(3'b011), .DQS_MODE(3'b011), .CDR_EN(2'b00)
        , .HS_IO_CLK_SEL(9'b111001000), .DLL_CODE_SEL(2'b00), .CDR_CLK_SEL(12'b000000000001)
        , .READ_MARGIN_TEST_EN(1'b0), .WRITE_MARGIN_TEST_EN(1'b1), .CDR_CLK_DIV(3'b000)
        , .DIV_CLK_SEL(2'b00), .HS_IO_CLK_PAUSE_EN(1'b1), .QDR_EN(1'b0)
        , .DYN_ODT_MODE(1'b0), .DIV_CLK_EN_SRC(2'b11), .RANK_2_MODE(1'b0)
         )  I_LANECTRL (.RX_DATA_VALID(RX_DATA_VALID), 
        .RX_BURST_DETECT(RX_BURST_DETECT), .RX_DELAY_LINE_OUT_OF_RANGE(
        RX_DELAY_LINE_OUT_OF_RANGE), .TX_DELAY_LINE_OUT_OF_RANGE(
        TX_DELAY_LINE_OUT_OF_RANGE), .CLK_OUT_R(CLK_OUT_R_0), 
        .A_OUT_RST_N(A_OUT_RST_N), .FAB_CLK(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .RESET(GND), .DDR_READ(GND), 
        .READ_CLK_SEL({GND, GND, GND}), .DELAY_LINE_SEL(GND), 
        .DELAY_LINE_LOAD(VCC), .DELAY_LINE_DIRECTION(GND), 
        .DELAY_LINE_MOVE(GND), .HS_IO_CLK_PAUSE(
        HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net), .DIV_CLK_EN_N(
        VCC), .RX_BIT_SLIP(GND), .CDR_CLK_A_SEL({GND, GND, GND, GND, 
        GND, GND, GND, GND}), .EYE_MONITOR_WIDTH_IN({GND, GND, GND}), 
        .ODT_EN(GND), .CODE_UPDATE(GND), .DQS(GND), .DQS_N(GND), 
        .HS_IO_CLK({GND, GND, GND, GND, 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0, 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90}), .DLL_CODE({GND, 
        GND, GND, GND, GND, GND, GND, GND}), .EYE_MONITOR_WIDTH_OUT({
        EYE_MONITOR_WIDTH_OUT[2], EYE_MONITOR_WIDTH_OUT[1], 
        EYE_MONITOR_WIDTH_OUT[0]}), .ODT_EN_SEL(ODT_EN_SEL_0), 
        .RX_DQS_90({RX_DQS_90_0[1], RX_DQS_90[0]}), .TX_DQS(TX_DQS), 
        .TX_DQS_270(TX_DQS_270), .FIFO_WR_PTR({FIFO_WR_PTR[2], 
        FIFO_WR_PTR[1], FIFO_WR_PTR[0]}), .FIFO_RD_PTR({FIFO_RD_PTR[2], 
        FIFO_RD_PTR[1], FIFO_RD_PTR[0]}), .CDR_CLK(CDR_CLK_0), 
        .CDR_NEXT_CLK(CDR_NEXT_CLK_0), .ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), .ODT_EN_OUT(ODT_EN_OUT_0), 
        .DDR_DO_READ(GND), .CDR_CLK_A_SEL_8(GND), .CDR_CLK_A_SEL_9(GND)
        , .CDR_CLK_A_SEL_10(GND), .CDR_CLK_B_SEL({GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .SWITCH(GND), 
        .CDR_CLR_NEXT_CLK_N(GND));
    PF_IOD_GENERIC_TX_C0_LANECTRL_ADDR_CMD_0_PF_LANECTRL_PAUSE_SYNC_1 
        I_LANECTRL_PAUSE_SYNC (.PF_IOD_TX_CCC_C0_0_TX_CLK_G(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net(
        HS_IO_CLK_PAUSE_SYNC_I_LANECTRL_PAUSE_SYNC_net), .OR2_PAUSE_Y(
        OR2_PAUSE_Y));
    VCC VCC_Z (.Y(VCC));
    CLKINT TX_DQS_inferred_clock_RNIIO99 (.A(TX_DQS), .Y(
        LANECTRL_ADDR_CMD_0_TX_DQS));
    CLKINT TX_DQS_270_inferred_clock_RNIA404 (.A(TX_DQS_270), .Y(
        LANECTRL_ADDR_CMD_0_TX_DQS_270));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_IOD_GENERIC_TX_C0(
       prbsgen_parallel_fab_0_prbs_out_msb_o_0,
       TXD_N,
       TXD,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX,
       TX_CLK_N,
       TX_CLK,
       PF_IOD_TX_CCC_C0_0_TX_CLK_G,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90,
       PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0,
       PLL_LOCK_c_i,
       N_81
    );
input  [7:0] prbsgen_parallel_fab_0_prbs_out_msb_o_0;
output [1:0] TXD_N;
output [1:0] TXD;
output [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
output TX_CLK_N;
output TX_CLK;
input  PF_IOD_TX_CCC_C0_0_TX_CLK_G;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90;
input  PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0;
input  PLL_LOCK_c_i;
input  N_81;

    wire OR2_PAUSE_Y, LANECTRL_ADDR_CMD_0_TX_SYNC_RST, 
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST, LANECTRL_ADDR_CMD_0_ARST_N, 
        LANECTRL_ADDR_CMD_0_TX_DQS_270, LANECTRL_ADDR_CMD_0_TX_DQS, 
        GND, VCC;
    
    PF_IOD_GENERIC_TX_C0_PF_IOD_TX_CLK_PF_IOD PF_IOD_TX_CLK (.TX_CLK(
        TX_CLK), .TX_CLK_N(TX_CLK_N), .LANECTRL_ADDR_CMD_0_TX_DQS_270(
        LANECTRL_ADDR_CMD_0_TX_DQS_270), .LANECTRL_ADDR_CMD_0_TX_DQS(
        LANECTRL_ADDR_CMD_0_TX_DQS), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90), 
        .LANECTRL_ADDR_CMD_0_TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), 
        .LANECTRL_ADDR_CMD_0_RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .LANECTRL_ADDR_CMD_0_ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .PF_IOD_TX_CCC_C0_0_TX_CLK_G(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G));
    OR2 OR2_PAUSE (.A(N_81), .B(PLL_LOCK_c_i), .Y(OR2_PAUSE_Y));
    PF_IOD_GENERIC_TX_C0_PF_IOD_TX_PF_IOD PF_IOD_TX (.TXD({TXD[1], 
        TXD[0]}), .TXD_N({TXD_N[1], TXD_N[0]}), 
        .prbsgen_parallel_fab_0_prbs_out_msb_o_0({
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[0]}), 
        .LANECTRL_ADDR_CMD_0_TX_DQS_270(LANECTRL_ADDR_CMD_0_TX_DQS_270)
        , .LANECTRL_ADDR_CMD_0_TX_DQS(LANECTRL_ADDR_CMD_0_TX_DQS), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0), 
        .LANECTRL_ADDR_CMD_0_TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), 
        .LANECTRL_ADDR_CMD_0_RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .LANECTRL_ADDR_CMD_0_ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .PF_IOD_TX_CCC_C0_0_TX_CLK_G(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G));
    PF_IOD_GENERIC_TX_C0_PF_IOD_CLK_TRAINING_PF_IOD 
        PF_IOD_CLK_TRAINING (
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX({
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]}), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0), 
        .LANECTRL_ADDR_CMD_0_TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), 
        .LANECTRL_ADDR_CMD_0_RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .LANECTRL_ADDR_CMD_0_ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), .PF_IOD_TX_CCC_C0_0_TX_CLK_G(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G));
    PF_IOD_GENERIC_TX_C0_LANECTRL_ADDR_CMD_0_PF_LANECTRL 
        LANECTRL_ADDR_CMD_0 (.OR2_PAUSE_Y(OR2_PAUSE_Y), 
        .LANECTRL_ADDR_CMD_0_TX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_TX_SYNC_RST), 
        .LANECTRL_ADDR_CMD_0_RX_SYNC_RST(
        LANECTRL_ADDR_CMD_0_RX_SYNC_RST), .LANECTRL_ADDR_CMD_0_ARST_N(
        LANECTRL_ADDR_CMD_0_ARST_N), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90), 
        .PF_IOD_TX_CCC_C0_0_TX_CLK_G(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .LANECTRL_ADDR_CMD_0_TX_DQS_270(LANECTRL_ADDR_CMD_0_TX_DQS_270)
        , .LANECTRL_ADDR_CMD_0_TX_DQS(LANECTRL_ADDR_CMD_0_TX_DQS));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module 
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_TRNG_Z1_1(
        
       BIT_ALGN_EYE_IN_c,
       EYE_MONITOR_EARLY_net_0_0,
       EYE_MONITOR_LATE_net_0_0,
       PLL_LOCK_0,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS,
       BIT_ALGN_DONE_c,
       BIT_ALGN_START_1_c,
       BIT_ALGN_OOR_c,
       BIT_ALGN_ERR_0_c,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD,
       debouncer_0_DB_OUT,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst
    );
input  [2:0] BIT_ALGN_EYE_IN_c;
input  EYE_MONITOR_EARLY_net_0_0;
input  EYE_MONITOR_LATE_net_0_0;
input  PLL_LOCK_0;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS;
output BIT_ALGN_DONE_c;
output BIT_ALGN_START_1_c;
input  BIT_ALGN_OOR_c;
output BIT_ALGN_ERR_0_c;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD;
input  debouncer_0_DB_OUT;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  RX_CLK_ALIGN_DONE_arst;

    wire [9:0] rst_cnt_Z;
    wire [8:0] rst_cnt_s;
    wire [127:0] late_flags_Z;
    wire [127:0] un10_early_flags;
    wire [127:0] late_flags_7_fast_Z;
    wire [50:49] late_flags_RNO_Z;
    wire [127:0] early_flags_Z;
    wire [127:0] early_flags_7_fast_Z;
    wire [50:49] early_flags_RNO_Z;
    wire [3:0] restart_edge_reg_Z;
    wire [2:0] restart_reg_Z;
    wire [6:0] tap_cnt_Z;
    wire [2:0] wait_cnt_Z;
    wire [2:0] wait_cnt_4_Z;
    wire [2:0] retrain_reg_Z;
    wire [1:1] cnt_Z;
    wire [1:1] cnt_RNO_Z;
    wire [6:0] tapcnt_final_Z;
    wire [6:0] tapcnt_final_13_1_Z;
    wire [6:0] no_early_no_late_val_st1_Z;
    wire [6:0] emflag_cnt_Z;
    wire [6:0] no_early_no_late_val_end2_Z;
    wire [4:0] bitalign_curr_state_Z;
    wire [4:0] bitalign_curr_state_34;
    wire [7:0] noearly_nolate_diff_nxt_8;
    wire [6:0] tapcnt_final_upd_Z;
    wire [1:0] tapcnt_final_upd_8_Z;
    wire [6:3] tapcnt_final_upd_8;
    wire [6:0] early_val_Z;
    wire [6:0] late_val_Z;
    wire [6:0] no_early_no_late_val_st2_Z;
    wire [7:0] early_late_diff_Z;
    wire [7:0] early_late_diff_8;
    wire [7:0] noearly_nolate_diff_start_7;
    wire [6:0] no_early_no_late_val_end1_Z;
    wire [7:0] timeout_cnt_Z;
    wire [7:0] timeout_cnt_s;
    wire [5:0] emflag_cnt_s;
    wire [6:6] emflag_cnt_s_Z;
    wire [9:9] rst_cnt_s_Z;
    wire [6:0] timeout_cnt_cry;
    wire [0:0] timeout_cnt_RNI9ABM_Y;
    wire [1:1] timeout_cnt_RNI8UO41_Y;
    wire [2:2] timeout_cnt_RNI8J6J1_Y;
    wire [3:3] timeout_cnt_RNI99K12_Y;
    wire [4:4] timeout_cnt_RNIB02G2_Y;
    wire [5:5] timeout_cnt_RNIEOFU2_Y;
    wire [7:7] timeout_cnt_RNO_FCO;
    wire [7:7] timeout_cnt_RNO_Y;
    wire [6:6] timeout_cnt_RNIIHTC3_Y;
    wire [0:0] emflag_cnt_cry_cy_S_0;
    wire [0:0] emflag_cnt_cry_cy_Y_0;
    wire [5:0] emflag_cnt_cry_Z;
    wire [5:0] emflag_cnt_cry_Y_0;
    wire [6:6] emflag_cnt_s_FCO;
    wire [6:6] emflag_cnt_s_Y;
    wire [0:0] un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_S;
    wire [0:0] un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_Y;
    wire [1:1] tapcnt_final_RNIOTM22_Y;
    wire [1:1] un1_tap_cnt_0_sqmuxa_14_0_Z;
    wire [2:2] tapcnt_final_RNI2SF33_Y;
    wire [3:3] tapcnt_final_RNIES844_Y;
    wire [4:4] tapcnt_final_RNISU155_Y;
    wire [6:6] tap_cnt_RNO_0_FCO;
    wire [6:6] tap_cnt_RNO_0_Y;
    wire [5:5] tapcnt_final_RNIC3R56_Y;
    wire [0:0] early_val_RNIT7HB3_S;
    wire [0:0] early_val_RNIT7HB3_Y;
    wire [0:0] early_val_RNI3L2D1_Z;
    wire [0:0] un1_no_early_no_late_val_end1_1_1_RNIHEIR_Z;
    wire [6:1] tapcnt_final_13_m1;
    wire [1:1] early_val_RNI0M2N6_Y;
    wire [1:1] early_val_RNI6O2D1_Z;
    wire [1:1] un1_no_early_no_late_val_end1_1_1_RNIJGIR_Z;
    wire [2:2] early_val_RNI9AK2A_Y;
    wire [2:2] early_val_RNI9R2D1_Z;
    wire [2:2] un1_no_early_no_late_val_end1_1_1_RNILIIR_Z;
    wire [3:3] early_val_RNIO46ED_Y;
    wire [3:3] early_val_RNICU2D1_Z;
    wire [3:3] un1_no_early_no_late_val_end1_1_1_RNINKIR_Z;
    wire [4:4] early_val_RNID5OPG_Y;
    wire [4:4] early_val_RNIF13D1_Z;
    wire [4:4] un1_no_early_no_late_val_end1_1_1_RNIPMIR_Z;
    wire [6:6] tapcnt_final_13_RNO_FCO;
    wire [6:6] tapcnt_final_13_RNO_Y;
    wire [5:5] early_val_RNI8CA5K_Y;
    wire [5:5] early_val_RNII43D1_Z;
    wire [5:5] un1_no_early_no_late_val_end1_1_1_RNIROIR_Z;
    wire [8:1] rst_cnt_cry_Z;
    wire [8:1] rst_cnt_cry_Y_0;
    wire [9:9] rst_cnt_s_FCO_0;
    wire [9:9] rst_cnt_s_Y_0;
    wire [6:1] tapcnt_final_13_Z;
    wire [96:0] un10_early_flags_1_Z;
    wire [69:0] un10_early_flags_2_Z;
    wire [100:0] un10_early_flags_2_0;
    wire [87:46] un10_early_flags_3_Z;
    wire [127:127] early_flags_dec;
    wire [6:0] un1_no_early_no_late_val_end1_1_1_Z;
    wire [6:0] un1_no_early_no_late_val_st1_1_1;
    wire [0:0] tapcnt_final_13_1_1_0_Z;
    wire [15:15] un10_early_flags_1_0;
    wire mv_dn_fg_0_sqmuxa_i_o2_Z, N_12_i, CO0_0, CO0_0_i, 
        un1_restart_trng_fg_5_Z, N_19_i, N_209, N_208, VCC, GND, 
        N_28_i, N_26_i, N_24_i, N_1497_i, N_1496_i, sig_re_train_Z, 
        Restart_trng_edge_det_Z, N_32_i, N_30_i, 
        no_early_no_late_val_st1_0_sqmuxa_i_Z, 
        no_early_no_late_val_end2_0_sqmuxa_i, un16_tapcnt_final_4, 
        un16_tapcnt_final_5, un16_tapcnt_final_6, un16_tapcnt_final_7, 
        tapcnt_final_upd_0_sqmuxa_i_Z, tapcnt_final_upd_8_cry_2_0_Y, 
        early_flags_0_sqmuxa_2_i, early_val_0_sqmuxa_1_i_Z, 
        un16_tapcnt_final_0, un16_tapcnt_final_1, un16_tapcnt_final_2, 
        un16_tapcnt_final_3, early_late_diff_0_sqmuxa_1_i, 
        un1_restart_trng_fg_8_Z, un10_tapcnt_final_4, 
        no_early_no_late_val_end1_0_sqmuxa_1_i, un10_tapcnt_final_5, 
        un10_tapcnt_final_6, un10_tapcnt_final_7, un10_tapcnt_final_0, 
        un10_tapcnt_final_1, un10_tapcnt_final_2, un10_tapcnt_final_3, 
        bit_align_start_Z, N_1439_i, bit_align_done_0_sqmuxa_3_i_Z, 
        bit_align_done_Z, bit_align_done_2_sqmuxa_Z, calc_done_Z, 
        N_1431_i, calc_done_0_sqmuxa_2_i_Z, rx_trng_done1_Z, N_1415_i, 
        rx_trng_done1_0_sqmuxa_i_Z, rx_BIT_ALGN_LOAD_9, 
        rx_BIT_ALGN_LOAD_0_sqmuxa_1_i_Z, late_last_set_Z, 
        early_late_diff_2_sqmuxa_Z, un1_restart_trng_fg_6_Z, 
        rx_BIT_ALGN_DIR_0_sqmuxa_2_i_Z, rx_BIT_ALGN_MOVE_2_sqmuxa_Z, 
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_i_Z, bit_align_dly_done_Z, 
        bit_align_dly_done_2_sqmuxa_Z, 
        bit_align_dly_done_0_sqmuxa_1_i_Z, rx_trng_done_Z, N_1403, 
        rx_trng_done_0_sqmuxa_i_Z, reset_dly_fg_Z, reset_dly_fg4_Z, 
        sig_rx_BIT_ALGN_CLR_FLGS_Z, sig_rx_BIT_ALGN_CLR_FLGS_11, 
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i_Z, rx_err_Z, N_1392, 
        rx_err_0_sqmuxa_1_i_Z, late_cur_set_Z, late_cur_set_2_sqmuxa_Z, 
        late_cur_set_0_sqmuxa_i_Z, early_cur_set_Z, 
        early_val_2_sqmuxa_Z, early_cur_set_0_sqmuxa_i_Z, 
        early_last_set_Z, early_last_set_2_sqmuxa_Z, 
        early_last_set_0_sqmuxa_i_Z, mv_up_fg_Z, 
        tapcnt_final_upd_2_sqmuxa_1, mv_up_fg_0_sqmuxa_i_0_Z, 
        mv_dn_fg_Z, tapcnt_final_upd_3_sqmuxa_1, 
        mv_dn_fg_0_sqmuxa_i_0_Z, timeout_cnte, emflag_cnte, 
        timeout_cnt_cry_cy, restart_trng_fg_RNIBNT7_S, 
        restart_trng_fg_RNIBNT7_Y, restart_trng_fg_i, 
        emflag_cnt_cry_cy, N_1456_1, un1_restart_trng_fg_9_0_443_0, 
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Z, 
        noearly_nolate_diff_nxt_8_cry_0_0_cy_S, 
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Y, 
        noearly_nolate_diff_nxt_8_cry_0, 
        noearly_nolate_diff_nxt_8_cry_0_0_Y, 
        noearly_nolate_diff_nxt_8_cry_1, 
        noearly_nolate_diff_nxt_8_cry_1_0_Y, 
        noearly_nolate_diff_nxt_8_cry_2, 
        noearly_nolate_diff_nxt_8_cry_2_0_Y, 
        noearly_nolate_diff_nxt_8_cry_3, 
        noearly_nolate_diff_nxt_8_cry_3_0_Y, 
        noearly_nolate_diff_nxt_8_cry_4, 
        noearly_nolate_diff_nxt_8_cry_4_0_Y, 
        noearly_nolate_diff_nxt_8_cry_5, 
        noearly_nolate_diff_nxt_8_cry_5_0_Y, 
        noearly_nolate_diff_nxt_8_s_7_FCO, 
        noearly_nolate_diff_nxt_8_s_7_Y, 
        noearly_nolate_diff_nxt_8_cry_6, 
        noearly_nolate_diff_nxt_8_cry_6_0_Y, 
        early_late_diff_8_cry_0_0_cy_Z, early_late_diff_8_cry_0_0_cy_S, 
        early_late_diff_8_cry_0_0_cy_Y, early_late_diff_8_cry_0, 
        early_late_diff_8_cry_0_0_Y, early_late_diff_8_cry_1, 
        early_late_diff_8_cry_1_0_Y, early_late_diff_8_cry_2, 
        early_late_diff_8_cry_2_0_Y, early_late_diff_8_cry_3, 
        early_late_diff_8_cry_3_0_Y, early_late_diff_8_cry_4, 
        early_late_diff_8_cry_4_0_Y, early_late_diff_8_cry_5, 
        early_late_diff_8_cry_5_0_Y, early_late_diff_8_s_7_FCO, 
        early_late_diff_8_s_7_Y, early_late_diff_8_cry_6, 
        early_late_diff_8_cry_6_0_Y, 
        noearly_nolate_diff_start_7_cry_0_0_cy_Z, 
        noearly_nolate_diff_start_7_cry_0_0_cy_S, 
        noearly_nolate_diff_start_7_cry_0_0_cy_Y, 
        noearly_nolate_diff_start_7_cry_0, 
        noearly_nolate_diff_start_7_cry_0_0_Y, 
        noearly_nolate_diff_start_7_cry_1, 
        noearly_nolate_diff_start_7_cry_1_0_Y, 
        noearly_nolate_diff_start_7_cry_2, 
        noearly_nolate_diff_start_7_cry_2_0_Y, 
        noearly_nolate_diff_start_7_cry_3, 
        noearly_nolate_diff_start_7_cry_3_0_Y, 
        noearly_nolate_diff_start_7_cry_4, 
        noearly_nolate_diff_start_7_cry_4_0_Y, 
        noearly_nolate_diff_start_7_cry_5, 
        noearly_nolate_diff_start_7_cry_5_0_Y, 
        noearly_nolate_diff_start_7_s_7_FCO, 
        noearly_nolate_diff_start_7_s_7_Y, 
        noearly_nolate_diff_start_7_cry_6, 
        noearly_nolate_diff_start_7_cry_6_0_Y, tap_cnt_17_i_m2_cry_0, 
        N_60, N_89, tap_cnt_17_i_m2_cry_1, N_79, tap_cnt_17_i_m2_cry_2, 
        N_78, tap_cnt_17_i_m2_cry_3, N_77, tap_cnt_17_i_m2_cry_4, N_76, 
        N_74, tap_cnt_17_i_m2_cry_5, N_75, tapcnt_final_13_m1_cry_0, 
        un1_bitalign_curr_state169_12_sn, tapcnt_final_13_m1_cry_1, 
        tapcnt_final_13_m1_cry_2, tapcnt_final_13_m1_cry_3, 
        tapcnt_final_13_m1_cry_4, tapcnt_final_3_sqmuxa_Z, 
        tapcnt_final_13_m1_axb_6_1, tapcnt_final_13_m1_cry_5, 
        tapcnt_final_upd_8_cry_2, tapcnt_final_upd_8_cry_2_0_S, N_100, 
        tapcnt_final_upd_8_cry_3, tapcnt_final_upd_8_cry_3_0_Y, 
        tapcnt_final_upd_8_cry_4, tapcnt_final_upd_8_cry_4_0_Y, 
        tapcnt_final_upd_8_s_6_FCO, tapcnt_final_upd_8_s_6_Y, 
        tapcnt_final_upd_8_cry_5, tapcnt_final_upd_8_cry_5_0_Y, 
        tapcnt_final27_cry_0_Z, tapcnt_final27_cry_0_S, 
        tapcnt_final27_cry_0_Y, tapcnt_final27_cry_1_Z, 
        tapcnt_final27_cry_1_S, tapcnt_final27_cry_1_Y, 
        tapcnt_final27_cry_2_Z, tapcnt_final27_cry_2_S, 
        tapcnt_final27_cry_2_Y, tapcnt_final27_cry_3_Z, 
        tapcnt_final27_cry_3_S, tapcnt_final27_cry_3_Y, 
        tapcnt_final27_cry_4_Z, tapcnt_final27_cry_4_S, 
        tapcnt_final27_cry_4_Y, tapcnt_final27_cry_5_Z, 
        tapcnt_final27_cry_5_S, tapcnt_final27_cry_5_Y, tapcnt_final27, 
        tapcnt_final27_cry_6_S, tapcnt_final27_cry_6_Y, 
        un16_tapcnt_final_cry_0_Z, un16_tapcnt_final_cry_0_S, 
        un16_tapcnt_final_cry_0_Y, un16_tapcnt_final_cry_1_Z, 
        un16_tapcnt_final_cry_1_S, un16_tapcnt_final_cry_1_Y, 
        un16_tapcnt_final_cry_2_Z, un16_tapcnt_final_cry_2_S, 
        un16_tapcnt_final_cry_2_Y, un16_tapcnt_final_cry_3_Z, 
        un16_tapcnt_final_cry_3_S, un16_tapcnt_final_cry_3_Y, 
        un16_tapcnt_final_cry_4_Z, un16_tapcnt_final_cry_4_S, 
        un16_tapcnt_final_cry_4_Y, un16_tapcnt_final_cry_5_Z, 
        un16_tapcnt_final_cry_5_S, un16_tapcnt_final_cry_5_Y, 
        un16_tapcnt_final_cry_6_Z, un16_tapcnt_final_cry_6_S, 
        un16_tapcnt_final_cry_6_Y, un16_tapcnt_final_cry_7_Z, 
        un16_tapcnt_final_cry_7_S, un16_tapcnt_final_cry_7_Y, 
        un1_early_late_diff_1_cry_0_Z, un1_early_late_diff_1_cry_0_S, 
        un1_early_late_diff_1_cry_0_Y, un1_early_late_diff_1_cry_1_Z, 
        un1_early_late_diff_1_cry_1_S, un1_early_late_diff_1_cry_1_Y, 
        un1_early_late_diff_1_cry_2_Z, un1_early_late_diff_1_cry_2_S, 
        un1_early_late_diff_1_cry_2_Y, un1_early_late_diff_1_cry_3_Z, 
        un1_early_late_diff_1_cry_3_S, un1_early_late_diff_1_cry_3_Y, 
        un1_early_late_diff_1_cry_4_Z, un1_early_late_diff_1_cry_4_S, 
        un1_early_late_diff_1_cry_4_Y, un1_early_late_diff_1_cry_5_Z, 
        un1_early_late_diff_1_cry_5_S, un1_early_late_diff_1_cry_5_Y, 
        un1_early_late_diff_1_cry_6_Z, un1_early_late_diff_1_cry_6_S, 
        un1_early_late_diff_1_cry_6_Y, un1_early_late_diff_1_cry_7_Z, 
        un1_early_late_diff_1_cry_7_S, un1_early_late_diff_1_cry_7_Y, 
        un10_tapcnt_final_cry_0_Z, un10_tapcnt_final_cry_0_S, 
        un10_tapcnt_final_cry_0_Y, un10_tapcnt_final_cry_1_Z, 
        un10_tapcnt_final_cry_1_S, un10_tapcnt_final_cry_1_Y, 
        un10_tapcnt_final_cry_2_Z, un10_tapcnt_final_cry_2_S, 
        un10_tapcnt_final_cry_2_Y, un10_tapcnt_final_cry_3_Z, 
        un10_tapcnt_final_cry_3_S, un10_tapcnt_final_cry_3_Y, 
        un10_tapcnt_final_cry_4_Z, un10_tapcnt_final_cry_4_S, 
        un10_tapcnt_final_cry_4_Y, un10_tapcnt_final_cry_5_Z, 
        un10_tapcnt_final_cry_5_S, un10_tapcnt_final_cry_5_Y, 
        un10_tapcnt_final_cry_6_Z, un10_tapcnt_final_cry_6_S, 
        un10_tapcnt_final_cry_6_Y, un10_tapcnt_final_cry_7_Z, 
        un10_tapcnt_final_cry_7_S, un10_tapcnt_final_cry_7_Y, 
        un1_early_late_diff_cry_0_Z, un1_early_late_diff_cry_0_S, 
        un1_early_late_diff_cry_0_Y, un1_early_late_diff_cry_1_Z, 
        un1_early_late_diff_cry_1_S, un1_early_late_diff_cry_1_Y, 
        un1_early_late_diff_cry_2_Z, un1_early_late_diff_cry_2_S, 
        un1_early_late_diff_cry_2_Y, un1_early_late_diff_cry_3_Z, 
        un1_early_late_diff_cry_3_S, un1_early_late_diff_cry_3_Y, 
        un1_early_late_diff_cry_4_Z, un1_early_late_diff_cry_4_S, 
        un1_early_late_diff_cry_4_Y, un1_early_late_diff_cry_5_Z, 
        un1_early_late_diff_cry_5_S, un1_early_late_diff_cry_5_Y, 
        un1_early_late_diff_cry_6_Z, un1_early_late_diff_cry_6_S, 
        un1_early_late_diff_cry_6_Y, un1_early_late_diff_cry_7_Z, 
        un1_early_late_diff_cry_7_S, un1_early_late_diff_cry_7_Y, 
        rst_cnt_s_715_FCO, rst_cnt_s_715_S, rst_cnt_s_715_Y, 
        late_flags_pmux_127_1_0_co1, late_flags_pmux_127_1_0_wmux_0_S, 
        late_flags_pmux, late_flags_pmux_126_1_1_wmux_10_Y, 
        late_flags_pmux_126_1_0_wmux_10_Y, late_flags_pmux_127_1_0_y0, 
        late_flags_pmux_127_1_0_co0, late_flags_pmux_127_1_0_wmux_S, 
        late_flags_pmux_63_1_1_wmux_10_Y, 
        late_flags_pmux_63_1_0_wmux_10_Y, early_flags_pmux_127_1_0_co1, 
        early_flags_pmux_127_1_0_wmux_0_S, early_flags_pmux, 
        early_flags_pmux_126_1_1_wmux_10_Y, 
        early_flags_pmux_126_1_0_wmux_10_Y, 
        early_flags_pmux_127_1_0_y0, early_flags_pmux_127_1_0_co0, 
        early_flags_pmux_127_1_0_wmux_S, 
        early_flags_pmux_63_1_1_wmux_10_Y, 
        early_flags_pmux_63_1_0_wmux_10_Y, m74_2_1_1_1_co1, 
        m74_2_1_1_wmux_0_S, N_75_0, N_29_i, N_116_mux, m74_2_1_1_1_y0, 
        m74_2_1_1_1_co0, m74_2_1_1_1_wmux_S, N_69, m74_1_0, 
        early_flags_pmux_63_1_1_co1_9, 
        early_flags_pmux_63_1_1_wmux_20_S, early_flags_pmux_63_1_1_y21, 
        early_flags_pmux_63_1_1_y3_0, early_flags_pmux_63_1_1_y1_0, 
        early_flags_pmux_63_1_1_y0_8, early_flags_pmux_63_1_1_co0_9, 
        early_flags_pmux_63_1_1_wmux_19_S, 
        early_flags_pmux_63_1_1_y5_0, early_flags_pmux_63_1_1_y7_0, 
        early_flags_pmux_63_1_1_co1_8, 
        early_flags_pmux_63_1_1_wmux_18_S, 
        early_flags_pmux_63_1_1_y0_7, early_flags_pmux_63_1_1_co0_8, 
        early_flags_pmux_63_1_1_wmux_17_S, 
        early_flags_pmux_63_1_1_co1_7, 
        early_flags_pmux_63_1_1_wmux_16_S, 
        early_flags_pmux_63_1_1_y0_6, early_flags_pmux_63_1_1_co0_7, 
        early_flags_pmux_63_1_1_wmux_15_S, 
        early_flags_pmux_63_1_1_co1_6, 
        early_flags_pmux_63_1_1_wmux_14_S, 
        early_flags_pmux_63_1_1_y0_5, early_flags_pmux_63_1_1_co0_6, 
        early_flags_pmux_63_1_1_wmux_13_S, 
        early_flags_pmux_63_1_1_co1_5, 
        early_flags_pmux_63_1_1_wmux_12_S, 
        early_flags_pmux_63_1_1_y0_4, early_flags_pmux_63_1_1_co0_5, 
        early_flags_pmux_63_1_1_wmux_11_S, 
        early_flags_pmux_63_1_1_co1_4, 
        early_flags_pmux_63_1_1_wmux_10_S, early_flags_pmux_63_1_1_y9, 
        early_flags_pmux_63_1_1_co0_4, 
        early_flags_pmux_63_1_1_wmux_9_S, 
        early_flags_pmux_63_1_1_wmux_9_Y, 
        early_flags_pmux_63_1_1_co1_3, 
        early_flags_pmux_63_1_1_wmux_8_S, early_flags_pmux_63_1_1_y3, 
        early_flags_pmux_63_1_1_y1, early_flags_pmux_63_1_1_y0_3, 
        early_flags_pmux_63_1_1_co0_3, 
        early_flags_pmux_63_1_1_wmux_7_S, early_flags_pmux_63_1_1_y5, 
        early_flags_pmux_63_1_1_y7, early_flags_pmux_63_1_1_co1_2, 
        early_flags_pmux_63_1_1_wmux_6_S, early_flags_pmux_63_1_1_y0_2, 
        early_flags_pmux_63_1_1_co0_2, 
        early_flags_pmux_63_1_1_wmux_5_S, 
        early_flags_pmux_63_1_1_co1_1, 
        early_flags_pmux_63_1_1_wmux_4_S, early_flags_pmux_63_1_1_y0_1, 
        early_flags_pmux_63_1_1_co0_1, 
        early_flags_pmux_63_1_1_wmux_3_S, 
        early_flags_pmux_63_1_1_co1_0, 
        early_flags_pmux_63_1_1_wmux_2_S, early_flags_pmux_63_1_1_y0_0, 
        early_flags_pmux_63_1_1_co0_0, 
        early_flags_pmux_63_1_1_wmux_1_S, early_flags_pmux_63_1_1_co1, 
        early_flags_pmux_63_1_1_wmux_0_S, early_flags_pmux_63_1_1_y0, 
        early_flags_pmux_63_1_1_co0, early_flags_pmux_63_1_1_wmux_S, 
        late_flags_pmux_126_1_1_co1_9, 
        late_flags_pmux_126_1_1_wmux_20_S, late_flags_pmux_126_1_1_y21, 
        late_flags_pmux_126_1_1_y3_0, late_flags_pmux_126_1_1_y1_0, 
        late_flags_pmux_126_1_1_y0_8, late_flags_pmux_126_1_1_co0_9, 
        late_flags_pmux_126_1_1_wmux_19_S, 
        late_flags_pmux_126_1_1_y5_0, late_flags_pmux_126_1_1_y7_0, 
        late_flags_pmux_126_1_1_co1_8, 
        late_flags_pmux_126_1_1_wmux_18_S, 
        late_flags_pmux_126_1_1_y0_7, late_flags_pmux_126_1_1_co0_8, 
        late_flags_pmux_126_1_1_wmux_17_S, 
        late_flags_pmux_126_1_1_co1_7, 
        late_flags_pmux_126_1_1_wmux_16_S, 
        late_flags_pmux_126_1_1_y0_6, late_flags_pmux_126_1_1_co0_7, 
        late_flags_pmux_126_1_1_wmux_15_S, 
        late_flags_pmux_126_1_1_co1_6, 
        late_flags_pmux_126_1_1_wmux_14_S, 
        late_flags_pmux_126_1_1_y0_5, late_flags_pmux_126_1_1_co0_6, 
        late_flags_pmux_126_1_1_wmux_13_S, 
        late_flags_pmux_126_1_1_co1_5, 
        late_flags_pmux_126_1_1_wmux_12_S, 
        late_flags_pmux_126_1_1_y0_4, late_flags_pmux_126_1_1_co0_5, 
        late_flags_pmux_126_1_1_wmux_11_S, 
        late_flags_pmux_126_1_1_co1_4, 
        late_flags_pmux_126_1_1_wmux_10_S, late_flags_pmux_126_1_1_y9, 
        late_flags_pmux_126_1_1_co0_4, 
        late_flags_pmux_126_1_1_wmux_9_S, 
        late_flags_pmux_126_1_1_wmux_9_Y, 
        late_flags_pmux_126_1_1_co1_3, 
        late_flags_pmux_126_1_1_wmux_8_S, late_flags_pmux_126_1_1_y3, 
        late_flags_pmux_126_1_1_y1, late_flags_pmux_126_1_1_y0_3, 
        late_flags_pmux_126_1_1_co0_3, 
        late_flags_pmux_126_1_1_wmux_7_S, late_flags_pmux_126_1_1_y5, 
        late_flags_pmux_126_1_1_y7, late_flags_pmux_126_1_1_co1_2, 
        late_flags_pmux_126_1_1_wmux_6_S, late_flags_pmux_126_1_1_y0_2, 
        late_flags_pmux_126_1_1_co0_2, 
        late_flags_pmux_126_1_1_wmux_5_S, 
        late_flags_pmux_126_1_1_co1_1, 
        late_flags_pmux_126_1_1_wmux_4_S, late_flags_pmux_126_1_1_y0_1, 
        late_flags_pmux_126_1_1_co0_1, 
        late_flags_pmux_126_1_1_wmux_3_S, 
        late_flags_pmux_126_1_1_co1_0, 
        late_flags_pmux_126_1_1_wmux_2_S, late_flags_pmux_126_1_1_y0_0, 
        late_flags_pmux_126_1_1_co0_0, 
        late_flags_pmux_126_1_1_wmux_1_S, late_flags_pmux_126_1_1_co1, 
        late_flags_pmux_126_1_1_wmux_0_S, late_flags_pmux_126_1_1_y0, 
        late_flags_pmux_126_1_1_co0, late_flags_pmux_126_1_1_wmux_S, 
        late_flags_pmux_63_1_0_co1_9, late_flags_pmux_63_1_0_wmux_20_S, 
        late_flags_pmux_63_1_0_0_y21, late_flags_pmux_63_1_0_y3_0, 
        late_flags_pmux_63_1_0_y1_0, late_flags_pmux_63_1_0_y0_8, 
        late_flags_pmux_63_1_0_co0_9, late_flags_pmux_63_1_0_wmux_19_S, 
        late_flags_pmux_63_1_0_y5_0, late_flags_pmux_63_1_0_y7_0, 
        late_flags_pmux_63_1_0_co1_8, late_flags_pmux_63_1_0_wmux_18_S, 
        late_flags_pmux_63_1_0_y0_7, late_flags_pmux_63_1_0_co0_8, 
        late_flags_pmux_63_1_0_wmux_17_S, late_flags_pmux_63_1_0_co1_7, 
        late_flags_pmux_63_1_0_wmux_16_S, late_flags_pmux_63_1_0_y0_6, 
        late_flags_pmux_63_1_0_co0_7, late_flags_pmux_63_1_0_wmux_15_S, 
        late_flags_pmux_63_1_0_co1_6, late_flags_pmux_63_1_0_wmux_14_S, 
        late_flags_pmux_63_1_0_y0_5, late_flags_pmux_63_1_0_co0_6, 
        late_flags_pmux_63_1_0_wmux_13_S, late_flags_pmux_63_1_0_co1_5, 
        late_flags_pmux_63_1_0_wmux_12_S, late_flags_pmux_63_1_0_y0_4, 
        late_flags_pmux_63_1_0_co0_5, late_flags_pmux_63_1_0_wmux_11_S, 
        late_flags_pmux_63_1_0_co1_4, late_flags_pmux_63_1_0_wmux_10_S, 
        late_flags_pmux_63_1_0_0_y9, late_flags_pmux_63_1_0_co0_4, 
        late_flags_pmux_63_1_0_wmux_9_S, 
        late_flags_pmux_63_1_0_wmux_9_Y, late_flags_pmux_63_1_0_co1_3, 
        late_flags_pmux_63_1_0_wmux_8_S, late_flags_pmux_63_1_0_0_y3, 
        late_flags_pmux_63_1_0_0_y1, late_flags_pmux_63_1_0_y0_3, 
        late_flags_pmux_63_1_0_co0_3, late_flags_pmux_63_1_0_wmux_7_S, 
        late_flags_pmux_63_1_0_0_y5, late_flags_pmux_63_1_0_0_y7, 
        late_flags_pmux_63_1_0_co1_2, late_flags_pmux_63_1_0_wmux_6_S, 
        late_flags_pmux_63_1_0_y0_2, late_flags_pmux_63_1_0_co0_2, 
        late_flags_pmux_63_1_0_wmux_5_S, late_flags_pmux_63_1_0_co1_1, 
        late_flags_pmux_63_1_0_wmux_4_S, late_flags_pmux_63_1_0_y0_1, 
        late_flags_pmux_63_1_0_co0_1, late_flags_pmux_63_1_0_wmux_3_S, 
        late_flags_pmux_63_1_0_co1_0, late_flags_pmux_63_1_0_wmux_2_S, 
        late_flags_pmux_63_1_0_y0_0, late_flags_pmux_63_1_0_co0_0, 
        late_flags_pmux_63_1_0_wmux_1_S, late_flags_pmux_63_1_0_0_co1, 
        late_flags_pmux_63_1_0_wmux_0_S, late_flags_pmux_63_1_0_0_y0, 
        late_flags_pmux_63_1_0_0_co0, late_flags_pmux_63_1_0_0_wmux_S, 
        early_flags_pmux_126_1_0_co1_9, 
        early_flags_pmux_126_1_0_wmux_20_S, 
        early_flags_pmux_126_1_0_0_y21, early_flags_pmux_126_1_0_y3_0, 
        early_flags_pmux_126_1_0_y1_0, early_flags_pmux_126_1_0_y0_8, 
        early_flags_pmux_126_1_0_co0_9, 
        early_flags_pmux_126_1_0_wmux_19_S, 
        early_flags_pmux_126_1_0_y5_0, early_flags_pmux_126_1_0_y7_0, 
        early_flags_pmux_126_1_0_co1_8, 
        early_flags_pmux_126_1_0_wmux_18_S, 
        early_flags_pmux_126_1_0_y0_7, early_flags_pmux_126_1_0_co0_8, 
        early_flags_pmux_126_1_0_wmux_17_S, 
        early_flags_pmux_126_1_0_co1_7, 
        early_flags_pmux_126_1_0_wmux_16_S, 
        early_flags_pmux_126_1_0_y0_6, early_flags_pmux_126_1_0_co0_7, 
        early_flags_pmux_126_1_0_wmux_15_S, 
        early_flags_pmux_126_1_0_co1_6, 
        early_flags_pmux_126_1_0_wmux_14_S, 
        early_flags_pmux_126_1_0_y0_5, early_flags_pmux_126_1_0_co0_6, 
        early_flags_pmux_126_1_0_wmux_13_S, 
        early_flags_pmux_126_1_0_co1_5, 
        early_flags_pmux_126_1_0_wmux_12_S, 
        early_flags_pmux_126_1_0_y0_4, early_flags_pmux_126_1_0_co0_5, 
        early_flags_pmux_126_1_0_wmux_11_S, 
        early_flags_pmux_126_1_0_co1_4, 
        early_flags_pmux_126_1_0_wmux_10_S, 
        early_flags_pmux_126_1_0_0_y9, early_flags_pmux_126_1_0_co0_4, 
        early_flags_pmux_126_1_0_wmux_9_S, 
        early_flags_pmux_126_1_0_wmux_9_Y, 
        early_flags_pmux_126_1_0_co1_3, 
        early_flags_pmux_126_1_0_wmux_8_S, 
        early_flags_pmux_126_1_0_0_y3, early_flags_pmux_126_1_0_0_y1, 
        early_flags_pmux_126_1_0_y0_3, early_flags_pmux_126_1_0_co0_3, 
        early_flags_pmux_126_1_0_wmux_7_S, 
        early_flags_pmux_126_1_0_0_y5, early_flags_pmux_126_1_0_0_y7, 
        early_flags_pmux_126_1_0_co1_2, 
        early_flags_pmux_126_1_0_wmux_6_S, 
        early_flags_pmux_126_1_0_y0_2, early_flags_pmux_126_1_0_co0_2, 
        early_flags_pmux_126_1_0_wmux_5_S, 
        early_flags_pmux_126_1_0_co1_1, 
        early_flags_pmux_126_1_0_wmux_4_S, 
        early_flags_pmux_126_1_0_y0_1, early_flags_pmux_126_1_0_co0_1, 
        early_flags_pmux_126_1_0_wmux_3_S, 
        early_flags_pmux_126_1_0_co1_0, 
        early_flags_pmux_126_1_0_wmux_2_S, 
        early_flags_pmux_126_1_0_y0_0, early_flags_pmux_126_1_0_co0_0, 
        early_flags_pmux_126_1_0_wmux_1_S, 
        early_flags_pmux_126_1_0_0_co1, 
        early_flags_pmux_126_1_0_wmux_0_S, 
        early_flags_pmux_126_1_0_0_y0, early_flags_pmux_126_1_0_0_co0, 
        early_flags_pmux_126_1_0_0_wmux_S, 
        early_flags_pmux_126_1_1_co1_9, 
        early_flags_pmux_126_1_1_wmux_20_S, 
        early_flags_pmux_126_1_1_y21, early_flags_pmux_126_1_1_y3_0, 
        early_flags_pmux_126_1_1_y1_0, early_flags_pmux_126_1_1_y0_8, 
        early_flags_pmux_126_1_1_co0_9, 
        early_flags_pmux_126_1_1_wmux_19_S, 
        early_flags_pmux_126_1_1_y5_0, early_flags_pmux_126_1_1_y7_0, 
        early_flags_pmux_126_1_1_co1_8, 
        early_flags_pmux_126_1_1_wmux_18_S, 
        early_flags_pmux_126_1_1_y0_7, early_flags_pmux_126_1_1_co0_8, 
        early_flags_pmux_126_1_1_wmux_17_S, 
        early_flags_pmux_126_1_1_co1_7, 
        early_flags_pmux_126_1_1_wmux_16_S, 
        early_flags_pmux_126_1_1_y0_6, early_flags_pmux_126_1_1_co0_7, 
        early_flags_pmux_126_1_1_wmux_15_S, 
        early_flags_pmux_126_1_1_co1_6, 
        early_flags_pmux_126_1_1_wmux_14_S, 
        early_flags_pmux_126_1_1_y0_5, early_flags_pmux_126_1_1_co0_6, 
        early_flags_pmux_126_1_1_wmux_13_S, 
        early_flags_pmux_126_1_1_co1_5, 
        early_flags_pmux_126_1_1_wmux_12_S, 
        early_flags_pmux_126_1_1_y0_4, early_flags_pmux_126_1_1_co0_5, 
        early_flags_pmux_126_1_1_wmux_11_S, 
        early_flags_pmux_126_1_1_co1_4, 
        early_flags_pmux_126_1_1_wmux_10_S, 
        early_flags_pmux_126_1_1_y9, early_flags_pmux_126_1_1_co0_4, 
        early_flags_pmux_126_1_1_wmux_9_S, 
        early_flags_pmux_126_1_1_wmux_9_Y, 
        early_flags_pmux_126_1_1_co1_3, 
        early_flags_pmux_126_1_1_wmux_8_S, early_flags_pmux_126_1_1_y3, 
        early_flags_pmux_126_1_1_y1, early_flags_pmux_126_1_1_y0_3, 
        early_flags_pmux_126_1_1_co0_3, 
        early_flags_pmux_126_1_1_wmux_7_S, early_flags_pmux_126_1_1_y5, 
        early_flags_pmux_126_1_1_y7, early_flags_pmux_126_1_1_co1_2, 
        early_flags_pmux_126_1_1_wmux_6_S, 
        early_flags_pmux_126_1_1_y0_2, early_flags_pmux_126_1_1_co0_2, 
        early_flags_pmux_126_1_1_wmux_5_S, 
        early_flags_pmux_126_1_1_co1_1, 
        early_flags_pmux_126_1_1_wmux_4_S, 
        early_flags_pmux_126_1_1_y0_1, early_flags_pmux_126_1_1_co0_1, 
        early_flags_pmux_126_1_1_wmux_3_S, 
        early_flags_pmux_126_1_1_co1_0, 
        early_flags_pmux_126_1_1_wmux_2_S, 
        early_flags_pmux_126_1_1_y0_0, early_flags_pmux_126_1_1_co0_0, 
        early_flags_pmux_126_1_1_wmux_1_S, 
        early_flags_pmux_126_1_1_co1, 
        early_flags_pmux_126_1_1_wmux_0_S, early_flags_pmux_126_1_1_y0, 
        early_flags_pmux_126_1_1_co0, early_flags_pmux_126_1_1_wmux_S, 
        early_flags_pmux_63_1_0_co1_9, 
        early_flags_pmux_63_1_0_wmux_20_S, 
        early_flags_pmux_63_1_0_0_y21, early_flags_pmux_63_1_0_y3_0, 
        early_flags_pmux_63_1_0_y1_0, early_flags_pmux_63_1_0_y0_8, 
        early_flags_pmux_63_1_0_co0_9, 
        early_flags_pmux_63_1_0_wmux_19_S, 
        early_flags_pmux_63_1_0_y5_0, early_flags_pmux_63_1_0_y7_0, 
        early_flags_pmux_63_1_0_co1_8, 
        early_flags_pmux_63_1_0_wmux_18_S, 
        early_flags_pmux_63_1_0_y0_7, early_flags_pmux_63_1_0_co0_8, 
        early_flags_pmux_63_1_0_wmux_17_S, 
        early_flags_pmux_63_1_0_co1_7, 
        early_flags_pmux_63_1_0_wmux_16_S, 
        early_flags_pmux_63_1_0_y0_6, early_flags_pmux_63_1_0_co0_7, 
        early_flags_pmux_63_1_0_wmux_15_S, 
        early_flags_pmux_63_1_0_co1_6, 
        early_flags_pmux_63_1_0_wmux_14_S, 
        early_flags_pmux_63_1_0_y0_5, early_flags_pmux_63_1_0_co0_6, 
        early_flags_pmux_63_1_0_wmux_13_S, 
        early_flags_pmux_63_1_0_co1_5, 
        early_flags_pmux_63_1_0_wmux_12_S, 
        early_flags_pmux_63_1_0_y0_4, early_flags_pmux_63_1_0_co0_5, 
        early_flags_pmux_63_1_0_wmux_11_S, 
        early_flags_pmux_63_1_0_co1_4, 
        early_flags_pmux_63_1_0_wmux_10_S, 
        early_flags_pmux_63_1_0_0_y9, early_flags_pmux_63_1_0_co0_4, 
        early_flags_pmux_63_1_0_wmux_9_S, 
        early_flags_pmux_63_1_0_wmux_9_Y, 
        early_flags_pmux_63_1_0_co1_3, 
        early_flags_pmux_63_1_0_wmux_8_S, early_flags_pmux_63_1_0_0_y3, 
        early_flags_pmux_63_1_0_0_y1, early_flags_pmux_63_1_0_y0_3, 
        early_flags_pmux_63_1_0_co0_3, 
        early_flags_pmux_63_1_0_wmux_7_S, early_flags_pmux_63_1_0_0_y5, 
        early_flags_pmux_63_1_0_0_y7, early_flags_pmux_63_1_0_co1_2, 
        early_flags_pmux_63_1_0_wmux_6_S, early_flags_pmux_63_1_0_y0_2, 
        early_flags_pmux_63_1_0_co0_2, 
        early_flags_pmux_63_1_0_wmux_5_S, 
        early_flags_pmux_63_1_0_co1_1, 
        early_flags_pmux_63_1_0_wmux_4_S, early_flags_pmux_63_1_0_y0_1, 
        early_flags_pmux_63_1_0_co0_1, 
        early_flags_pmux_63_1_0_wmux_3_S, 
        early_flags_pmux_63_1_0_co1_0, 
        early_flags_pmux_63_1_0_wmux_2_S, early_flags_pmux_63_1_0_y0_0, 
        early_flags_pmux_63_1_0_co0_0, 
        early_flags_pmux_63_1_0_wmux_1_S, 
        early_flags_pmux_63_1_0_0_co1, 
        early_flags_pmux_63_1_0_wmux_0_S, early_flags_pmux_63_1_0_0_y0, 
        early_flags_pmux_63_1_0_0_co0, 
        early_flags_pmux_63_1_0_0_wmux_S, late_flags_pmux_63_1_1_co1_9, 
        late_flags_pmux_63_1_1_wmux_20_S, late_flags_pmux_63_1_1_y21, 
        late_flags_pmux_63_1_1_y3_0, late_flags_pmux_63_1_1_y1_0, 
        late_flags_pmux_63_1_1_y0_8, late_flags_pmux_63_1_1_co0_9, 
        late_flags_pmux_63_1_1_wmux_19_S, late_flags_pmux_63_1_1_y5_0, 
        late_flags_pmux_63_1_1_y7_0, late_flags_pmux_63_1_1_co1_8, 
        late_flags_pmux_63_1_1_wmux_18_S, late_flags_pmux_63_1_1_y0_7, 
        late_flags_pmux_63_1_1_co0_8, late_flags_pmux_63_1_1_wmux_17_S, 
        late_flags_pmux_63_1_1_co1_7, late_flags_pmux_63_1_1_wmux_16_S, 
        late_flags_pmux_63_1_1_y0_6, late_flags_pmux_63_1_1_co0_7, 
        late_flags_pmux_63_1_1_wmux_15_S, late_flags_pmux_63_1_1_co1_6, 
        late_flags_pmux_63_1_1_wmux_14_S, late_flags_pmux_63_1_1_y0_5, 
        late_flags_pmux_63_1_1_co0_6, late_flags_pmux_63_1_1_wmux_13_S, 
        late_flags_pmux_63_1_1_co1_5, late_flags_pmux_63_1_1_wmux_12_S, 
        late_flags_pmux_63_1_1_y0_4, late_flags_pmux_63_1_1_co0_5, 
        late_flags_pmux_63_1_1_wmux_11_S, late_flags_pmux_63_1_1_co1_4, 
        late_flags_pmux_63_1_1_wmux_10_S, late_flags_pmux_63_1_1_y9, 
        late_flags_pmux_63_1_1_co0_4, late_flags_pmux_63_1_1_wmux_9_S, 
        late_flags_pmux_63_1_1_wmux_9_Y, late_flags_pmux_63_1_1_co1_3, 
        late_flags_pmux_63_1_1_wmux_8_S, late_flags_pmux_63_1_1_y3, 
        late_flags_pmux_63_1_1_y1, late_flags_pmux_63_1_1_y0_3, 
        late_flags_pmux_63_1_1_co0_3, late_flags_pmux_63_1_1_wmux_7_S, 
        late_flags_pmux_63_1_1_y5, late_flags_pmux_63_1_1_y7, 
        late_flags_pmux_63_1_1_co1_2, late_flags_pmux_63_1_1_wmux_6_S, 
        late_flags_pmux_63_1_1_y0_2, late_flags_pmux_63_1_1_co0_2, 
        late_flags_pmux_63_1_1_wmux_5_S, late_flags_pmux_63_1_1_co1_1, 
        late_flags_pmux_63_1_1_wmux_4_S, late_flags_pmux_63_1_1_y0_1, 
        late_flags_pmux_63_1_1_co0_1, late_flags_pmux_63_1_1_wmux_3_S, 
        late_flags_pmux_63_1_1_co1_0, late_flags_pmux_63_1_1_wmux_2_S, 
        late_flags_pmux_63_1_1_y0_0, late_flags_pmux_63_1_1_co0_0, 
        late_flags_pmux_63_1_1_wmux_1_S, late_flags_pmux_63_1_1_co1, 
        late_flags_pmux_63_1_1_wmux_0_S, late_flags_pmux_63_1_1_y0, 
        late_flags_pmux_63_1_1_co0, late_flags_pmux_63_1_1_wmux_S, 
        late_flags_pmux_126_1_0_co1_9, 
        late_flags_pmux_126_1_0_wmux_20_S, 
        late_flags_pmux_126_1_0_0_y21, late_flags_pmux_126_1_0_y3_0, 
        late_flags_pmux_126_1_0_y1_0, late_flags_pmux_126_1_0_y0_8, 
        late_flags_pmux_126_1_0_co0_9, 
        late_flags_pmux_126_1_0_wmux_19_S, 
        late_flags_pmux_126_1_0_y5_0, late_flags_pmux_126_1_0_y7_0, 
        late_flags_pmux_126_1_0_co1_8, 
        late_flags_pmux_126_1_0_wmux_18_S, 
        late_flags_pmux_126_1_0_y0_7, late_flags_pmux_126_1_0_co0_8, 
        late_flags_pmux_126_1_0_wmux_17_S, 
        late_flags_pmux_126_1_0_co1_7, 
        late_flags_pmux_126_1_0_wmux_16_S, 
        late_flags_pmux_126_1_0_y0_6, late_flags_pmux_126_1_0_co0_7, 
        late_flags_pmux_126_1_0_wmux_15_S, 
        late_flags_pmux_126_1_0_co1_6, 
        late_flags_pmux_126_1_0_wmux_14_S, 
        late_flags_pmux_126_1_0_y0_5, late_flags_pmux_126_1_0_co0_6, 
        late_flags_pmux_126_1_0_wmux_13_S, 
        late_flags_pmux_126_1_0_co1_5, 
        late_flags_pmux_126_1_0_wmux_12_S, 
        late_flags_pmux_126_1_0_y0_4, late_flags_pmux_126_1_0_co0_5, 
        late_flags_pmux_126_1_0_wmux_11_S, 
        late_flags_pmux_126_1_0_co1_4, 
        late_flags_pmux_126_1_0_wmux_10_S, 
        late_flags_pmux_126_1_0_0_y9, late_flags_pmux_126_1_0_co0_4, 
        late_flags_pmux_126_1_0_wmux_9_S, 
        late_flags_pmux_126_1_0_wmux_9_Y, 
        late_flags_pmux_126_1_0_co1_3, 
        late_flags_pmux_126_1_0_wmux_8_S, late_flags_pmux_126_1_0_0_y3, 
        late_flags_pmux_126_1_0_0_y1, late_flags_pmux_126_1_0_y0_3, 
        late_flags_pmux_126_1_0_co0_3, 
        late_flags_pmux_126_1_0_wmux_7_S, late_flags_pmux_126_1_0_0_y5, 
        late_flags_pmux_126_1_0_0_y7, late_flags_pmux_126_1_0_co1_2, 
        late_flags_pmux_126_1_0_wmux_6_S, late_flags_pmux_126_1_0_y0_2, 
        late_flags_pmux_126_1_0_co0_2, 
        late_flags_pmux_126_1_0_wmux_5_S, 
        late_flags_pmux_126_1_0_co1_1, 
        late_flags_pmux_126_1_0_wmux_4_S, late_flags_pmux_126_1_0_y0_1, 
        late_flags_pmux_126_1_0_co0_1, 
        late_flags_pmux_126_1_0_wmux_3_S, 
        late_flags_pmux_126_1_0_co1_0, 
        late_flags_pmux_126_1_0_wmux_2_S, late_flags_pmux_126_1_0_y0_0, 
        late_flags_pmux_126_1_0_co0_0, 
        late_flags_pmux_126_1_0_wmux_1_S, 
        late_flags_pmux_126_1_0_0_co1, 
        late_flags_pmux_126_1_0_wmux_0_S, late_flags_pmux_126_1_0_0_y0, 
        late_flags_pmux_126_1_0_0_co0, 
        late_flags_pmux_126_1_0_0_wmux_S, un1_bitalign_curr_state_12_Z, 
        un1_restart_trng_fg_10_sn, bitalign_curr_state12_Z, 
        bitalign_curr_state148_Z, bitalign_curr_state_1_sqmuxa_4_Z, 
        un1_tap_cnt_0_sqmuxa_6_0, bitalign_curr_state154_Z, 
        bitalign_curr_state164_Z, bitalign_curr_state41_Z, 
        calc_done_0_sqmuxa_Z, un1_bitalign_curr_state148_9_0_Z, un34, 
        calc_done25_Z, un1_noearly_nolate_diff_start_valid_Z, 
        calc_done27_Z, bitalign_curr_state160_Z, emflag_cnt_0_sqmuxa, 
        bitalign_curr_state159_Z, un1_early_last_set_1_sqmuxa_1_1_tz_Z, 
        bitalign_curr_state162_Z, un1_calc_done25_5_Z, 
        un1_early_late_diff_valid_Z, un10_early_flags_47_0_Z, 
        un10_early_flags_30_0_Z, N_20, late_last_set15_Z, N_94, N_60_0, 
        N_98, bitalign_curr_state148_2_Z, N_40, m40_1_1, 
        un1_restart_trng_fg_10_sn_1, early_last_set_1_sqmuxa_1_3_Z, 
        early_val_0_sqmuxa_1_0_Z, tap_cnt_0_sqmuxa_1_Z, N_100_0, 
        m101_1_1, N_102, bitalign_curr_state161_2_Z, N_92, m91_1, 
        m91_1_0, un1_retrain_adj_tap_i, m82_1_0, m82_1_1, N_83, 
        bitalign_curr_state89_Z, N_63, sig_rx_BIT_ALGN_CLR_FLGS14_Z, 
        m64_1_1, N_65, N_117_mux_1, m23_1_2, N_124_mux, m37_1_1, m37, 
        i12_mux_0, N_35, m7_1_1, N_8, tapcnt_final_2_sqmuxa_Z, m86_1, 
        m85_1, N_76_0, m67_1, m66_1, N_51, N_119_mux, m55_0, 
        tapcnt_final_13_m0s2_Z, un1_tapcnt_final_0_sqmuxa_Z, N_15, 
        m50_1_1, N_47, N_50, N_9, N_11, early_cur_set_0_sqmuxa_1_Z, 
        tapcnt_final_5_sqmuxa, rx_err_1_sqmuxa_Z, 
        calc_done_4_sqmuxa_0_Z, un1_bitalign_curr_state_0_sqmuxa_9_4_Z, 
        un1_bitalign_curr_state_0_sqmuxa_9_i, calc_done25_248_Z, 
        calc_done25_253_Z, calc_done25_249_Z, calc_done25_234_Z, 
        calc_done25_235_Z, calc_done25_251_Z, calc_done25_244_Z, 
        un1_bitalign_curr_state148_5_4_Z, 
        un1_bitalign_curr_state148_5_Z, calc_done25_160_Z, 
        calc_done25_161_Z, calc_done25_233_Z, calc_done25_209_Z, 
        un34lto7_3_Z, tap_cnt_0_sqmuxa_0_Z, rx_BIT_ALGN_ERR_3_Z, 
        reset_dly_fg4_4_Z, early_late_diff_0_sqmuxa_1_0_Z, 
        tap_cnt_0_sqmuxa_2_0, un1_bitalign_curr_state_1_sqmuxa_2_i_0, 
        N_63_0, rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z, N_82, N_1498, N_1499, 
        N_1416, i22_mux_1, un1_rx_BIT_ALGN_START, 
        bitalign_curr_state152_1_Z, tapcnt_final_upd_1_sqmuxa, 
        un1_sig_re_train_Z, bitalign_curr_state163_2, 
        un1_bitalign_curr_state_15_1_Z, bitalign_curr_state155_1_Z, 
        bitalign_curr_state159_2_Z, un1_early_flags_pmux_1_Z, 
        calc_done25_191_Z, calc_done25_190_Z, calc_done25_189_Z, 
        calc_done25_188_Z, calc_done25_187_Z, calc_done25_186_Z, 
        calc_done25_185_Z, calc_done25_184_Z, calc_done25_183_Z, 
        calc_done25_182_Z, calc_done25_181_Z, calc_done25_180_Z, 
        calc_done25_179_Z, calc_done25_178_Z, calc_done25_177_Z, 
        calc_done25_176_Z, calc_done25_175_Z, calc_done25_174_Z, 
        calc_done25_173_Z, calc_done25_172_Z, calc_done25_171_Z, 
        calc_done25_170_Z, calc_done25_169_Z, calc_done25_168_Z, 
        calc_done25_167_Z, calc_done25_166_Z, calc_done25_165_Z, 
        calc_done25_164_Z, calc_done25_163_Z, calc_done25_162_Z, 
        calc_done25_159_Z, calc_done25_158_Z, calc_done25_157_Z, 
        calc_done25_156_Z, calc_done25_155_Z, calc_done25_154_Z, 
        calc_done25_153_Z, calc_done25_152_Z, calc_done25_151_Z, 
        calc_done25_150_Z, calc_done25_149_Z, calc_done25_148_Z, 
        calc_done25_147_Z, calc_done25_146_Z, calc_done25_145_Z, 
        calc_done25_144_Z, calc_done25_143_Z, calc_done25_142_Z, 
        calc_done25_141_Z, calc_done25_140_Z, calc_done25_139_Z, 
        calc_done25_138_Z, calc_done25_137_Z, calc_done25_136_Z, 
        calc_done25_135_Z, calc_done25_134_Z, calc_done25_133_Z, 
        calc_done25_132_Z, calc_done25_131_Z, calc_done25_130_Z, 
        calc_done25_129_Z, calc_done25_128_Z, 
        bitalign_curr_state_2_sqmuxa_4_0_0_Z, 
        un2_noearly_nolate_diff_start_validlto7_2_Z, 
        un2_noearly_nolate_diff_nxt_validlto7_2_Z, 
        early_flags_dec_127_4_Z, un2_early_late_diff_validlto7_2_Z, 
        rx_BIT_ALGN_MOVE_0_sqmuxa_0_Z, un34lto7_4_Z, 
        tap_cnt_0_sqmuxa_1_0_Z, rx_BIT_ALGN_ERR_4_Z, reset_dly_fg4_6_Z, 
        un1_early_flags_1_sqmuxa_i, bitalign_curr_state_0_sqmuxa_10, 
        bitalign_curr_state61, N_114_mux, 
        un2_noearly_nolate_diff_nxt_validlt3, bitalign_curr_state13, 
        un1_bitalign_curr_state151_Z, bitalign_curr_state152_3_Z, 
        bitalign_curr_state154_3_Z, 
        un2_noearly_nolate_diff_start_validlt3, N_31, 
        un1_bitalign_curr_state_16_1_Z, bitalign_curr_state12_0, 
        reset_dly_fg4_8_Z, bitalign_curr_state161_Z, 
        bit_align_dly_done_0_sqmuxa_Z, bitalign_curr_state155_Z, 
        bitalign_curr_state_0_sqmuxa_8_Z, bitalign_curr_state153_Z, 
        bitalign_curr_state156_Z, bitalign_curr_state163_Z, N_108, 
        bitalign_curr_state149_Z, tapcnt_final_1_sqmuxa_2_Z, N_61, 
        un1_bitalign_curr_state152_Z, un1_restart_trng_fg_Z, 
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z, 
        un1_bitalign_curr_state_1_sqmuxa_6_i_0, 
        un2_early_late_diff_validlt7, un1_calc_done25_7_i, 
        bitalign_curr_state61_0, bitalign_curr_state61_1_Z, 
        bitalign_curr_state61_4_Z, bitalign_curr_state61_5_Z, 
        bitalign_curr_state61_6_Z, bitalign_curr_state61_3_Z, 
        bitalign_curr_state61_2_Z, un1_bitalign_curr_state_15_0_Z, 
        calc_done25_239_Z, calc_done25_238_Z, calc_done25_237_Z, 
        calc_done25_236_Z, calc_done25_231_Z, calc_done25_230_Z, 
        calc_done25_229_Z, calc_done25_228_Z, calc_done25_227_Z, 
        calc_done25_226_Z, calc_done25_225_Z, calc_done25_224_Z, 
        un1_bitalign_curr_state148_2_Z, rx_BIT_ALGN_LOAD_0_sqmuxa_Z, 
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_Z, 
        un1_bitalign_curr_state148_3_Z, early_flags_0_sqmuxa_1_Z, 
        early_flags_1_sqmuxa_1_Z, bit_align_done_0_sqmuxa_2_Z, N_52, 
        rx_trng_done_1_sqmuxa_Z, early_flags_0_sqmuxa_Z, 
        early_flags_1_sqmuxa_Z, CO1, un1_tapcnt_final_Z, 
        rx_BIT_ALGN_DIR_1_sqmuxa_Z, un1_rx_BIT_ALGN_LOAD_0_sqmuxa_i_0, 
        N_14, timeout_cntlde_0, un1_bitalign_curr_state148_8_0_Z, 
        un1_bitalign_curr_state148_4_1_Z, 
        bitalign_curr_state_0_sqmuxa_9_Z, 
        bit_align_done_0_sqmuxa_3_1_Z, early_late_diff_0_sqmuxa_Z, 
        un1_bitalign_curr_state_13_1_Z, un1_early_flags_1_sqmuxa_1_Z, 
        tapcnt_final_upd_3_sqmuxa_Z, 
        un1_noearly_nolate_diff_nxt_valid_Z, 
        bitalign_curr_state61_NE_4_Z, emflag_cntlde_1, 
        un1_bitalign_curr_state_0_sqmuxa_9_1_Z, 
        un1_restart_trng_fg_10_0_Z, rx_BIT_ALGN_MOVE_0_sqmuxa_2_1_Z, 
        un1_bitalign_curr_state_14_1_Z, 
        un1_bitalign_curr_state_2_sqmuxa_Z, i22_mux, 
        tapcnt_final_upd_2_sqmuxa, emflag_cnt_1_sqmuxa_1_Z, N_130_mux, 
        un1_bitalign_curr_state148_8_2_Z, 
        un1_bitalign_curr_state_15_3_Z, emflag_cntlde_4, 
        un1_bitalign_curr_state148_9_2_Z, calc_done26_Z, calc_done28_Z, 
        un1_bitalign_curr_state_0_sqmuxa_9_2_Z;
    
    SLE \cnt[0]  (.D(CO0_0_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(CO0_0));
    SLE \early_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[4]));
    CFG3 #( .INIT(8'h40) )  rx_BIT_ALGN_MOVE_0_sqmuxa_0 (.A(
        bitalign_curr_state_Z[0]), .B(tap_cnt_0_sqmuxa_2_0), .C(
        bitalign_curr_state_Z[1]), .Y(rx_BIT_ALGN_MOVE_0_sqmuxa_0_Z));
    SLE \late_flags[59]  (.D(late_flags_7_fast_Z[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[59]));
    SLE \early_flags[93]  (.D(early_flags_7_fast_Z[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[93]));
    CFG4 #( .INIT(16'h00CA) )  \bitalign_curr_state_34_4_0_.m112  (.A(
        i22_mux), .B(N_130_mux), .C(bitalign_curr_state_Z[4]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[4]));
    CFG3 #( .INIT(8'h04) )  \bitalign_curr_state_34_4_0_.m103  (.A(
        un1_bitalign_curr_state_0_sqmuxa_9_i), .B(N_102), .C(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[46]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[46]), .C(
        un10_early_flags[46]), .Y(late_flags_7_fast_Z[46]));
    SLE \late_flags[38]  (.D(late_flags_7_fast_Z[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[38]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[27]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[27]), .C(
        un10_early_flags[27]), .Y(early_flags_7_fast_Z[27]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[125]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[125]), .C(
        un10_early_flags[125]), .Y(early_flags_7_fast_Z[125]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_3 (.A(
        un10_early_flags_2_0[0]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[3]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[87]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[87]), .C(
        un10_early_flags[87]), .Y(early_flags_7_fast_Z[87]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[124]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[124]), .C(
        un10_early_flags[124]), .Y(early_flags_7_fast_Z[124]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[61]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[61]), .C(
        un10_early_flags[61]), .Y(late_flags_7_fast_Z[61]));
    SLE \early_flags[127]  (.D(early_flags_7_fast_Z[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[127]));
    CFG4 #( .INIT(16'h0008) )  bitalign_curr_state12 (.A(
        reset_dly_fg_Z), .B(bitalign_curr_state12_0), .C(
        BIT_ALGN_ERR_0_c), .D(rx_trng_done_Z), .Y(
        bitalign_curr_state12_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_30 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[0]), .D(un10_early_flags_30_0_Z), .Y(
        un10_early_flags[30]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_10 (.A(
        late_flags_pmux_63_1_0_0_y21), .B(late_flags_pmux_63_1_0_0_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_63_1_0_co0_4), .S(
        late_flags_pmux_63_1_0_wmux_10_S), .Y(
        late_flags_pmux_63_1_0_wmux_10_Y), .FCO(
        late_flags_pmux_63_1_0_co1_4));
    SLE \late_flags[95]  (.D(late_flags_7_fast_Z[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[95]));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_82 (.A(tap_cnt_Z[5]), 
        .B(N_1499), .C(un10_early_flags_2_Z[0]), .D(
        un10_early_flags_1_Z[64]), .Y(un10_early_flags[82]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[14]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[14]), .C(
        un10_early_flags[14]), .Y(late_flags_7_fast_Z[14]));
    SLE \late_flags[24]  (.D(late_flags_7_fast_Z[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[24]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_16 (.A(
        early_flags_pmux_126_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[45]), .D(early_flags_Z[109]), .FCI(
        early_flags_pmux_126_1_1_co0_7), .S(
        early_flags_pmux_126_1_1_wmux_16_S), .Y(
        early_flags_pmux_126_1_1_y5_0), .FCO(
        early_flags_pmux_126_1_1_co1_7));
    CFG2 #( .INIT(4'hB) )  rx_trng_done1_1_sqmuxa_i (.A(N_61), .B(
        bitalign_curr_state148_Z), .Y(N_52));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[82]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[82]), .C(
        un10_early_flags[82]), .Y(late_flags_7_fast_Z[82]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI3L2D1[0]  (.A(early_val_Z[0])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[0]), .Y(
        early_val_RNI3L2D1_Z[0]));
    SLE \late_flags[6]  (.D(late_flags_7_fast_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[67]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[67]), .C(
        un10_early_flags[67]), .Y(early_flags_7_fast_Z[67]));
    CFG3 #( .INIT(8'h01) )  bitalign_curr_state41 (.A(wait_cnt_Z[2]), 
        .B(wait_cnt_Z[1]), .C(wait_cnt_Z[0]), .Y(
        bitalign_curr_state41_Z));
    SLE \noearly_nolate_diff_start[7]  (.D(
        noearly_nolate_diff_start_7[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_7));
    CFG4 #( .INIT(16'h0C5C) )  \bitalign_curr_state_34_4_0_.m62  (.A(
        N_35), .B(N_60_0), .C(bitalign_curr_state_Z[0]), .D(
        early_flags_dec[127]), .Y(N_63));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_2 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[0]), .D(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[2]));
    SLE rx_trng_done1 (.D(N_1415_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_trng_done1_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_trng_done1_Z));
    CFG3 #( .INIT(8'hFB) )  bit_align_dly_done_0_sqmuxa_1_i (.A(
        tap_cnt_0_sqmuxa_1_Z), .B(bit_align_done_0_sqmuxa_3_1_Z), .C(
        bitalign_curr_state_0_sqmuxa_9_Z), .Y(
        bit_align_dly_done_0_sqmuxa_1_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[92]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[92]), .C(
        un10_early_flags[92]), .Y(early_flags_7_fast_Z[92]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_140 (.A(late_flags_Z[71]), 
        .B(late_flags_Z[70]), .C(late_flags_Z[69]), .D(
        late_flags_Z[68]), .Y(calc_done25_140_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_20 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[16]), .C(
        un10_early_flags_1_Z[20]), .Y(un10_early_flags[20]));
    SLE \late_flags[69]  (.D(late_flags_7_fast_Z[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[69]));
    CFG4 #( .INIT(16'h5540) )  early_val_2_sqmuxa (.A(
        restart_trng_fg_i), .B(un1_early_last_set_1_sqmuxa_1_1_tz_Z), 
        .C(early_flags_pmux), .D(early_last_set_1_sqmuxa_1_3_Z), .Y(
        early_val_2_sqmuxa_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_0 (.A(
        late_flags_pmux_63_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[34]), .D(late_flags_Z[98]), .FCI(
        late_flags_pmux_63_1_0_0_co0), .S(
        late_flags_pmux_63_1_0_wmux_0_S), .Y(
        late_flags_pmux_63_1_0_0_y1), .FCO(
        late_flags_pmux_63_1_0_0_co1));
    SLE rx_BIT_ALGN_LOAD (.D(rx_BIT_ALGN_LOAD_9), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_BIT_ALGN_LOAD_0_sqmuxa_1_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD));
    CFG4 #( .INIT(16'h8000) )  calc_done25_231 (.A(calc_done25_159_Z), 
        .B(calc_done25_158_Z), .C(calc_done25_157_Z), .D(
        calc_done25_156_Z), .Y(calc_done25_231_Z));
    SLE \late_flags[125]  (.D(late_flags_7_fast_Z[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[125]));
    SLE \early_late_diff[1]  (.D(early_late_diff_8[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[1]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNIB02G2[4]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[4]), .D(GND), .FCI(
        timeout_cnt_cry[3]), .S(timeout_cnt_s[4]), .Y(
        timeout_cnt_RNIB02G2_Y[4]), .FCO(timeout_cnt_cry[4]));
    CFG4 #( .INIT(16'h0010) )  bitalign_curr_state153 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        N_1456_1), .D(bitalign_curr_state_Z[1]), .Y(
        bitalign_curr_state153_Z));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_6 (.A(
        un10_tapcnt_final_6), .B(un16_tapcnt_final_6), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_5_Z), .S(
        un10_tapcnt_final_cry_6_S), .Y(un10_tapcnt_final_cry_6_Y), 
        .FCO(un10_tapcnt_final_cry_6_Z));
    SLE \late_flags[74]  (.D(late_flags_7_fast_Z[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[74]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_94 (.A(tap_cnt_Z[5]), 
        .B(un10_early_flags_1_Z[6]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[64]), .Y(un10_early_flags[94]));
    SLE \early_flags[34]  (.D(early_flags_7_fast_Z[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[34]));
    CFG4 #( .INIT(16'hF800) )  un1_noearly_nolate_diff_nxt_valid (.A(
        un16_tapcnt_final_3), .B(un2_noearly_nolate_diff_nxt_validlt3), 
        .C(un2_noearly_nolate_diff_nxt_validlto7_2_Z), .D(
        un1_early_late_diff_1_cry_7_Z), .Y(
        un1_noearly_nolate_diff_nxt_valid_Z));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIT7HB3[0]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIHEIR_Z[0]), .B(
        early_val_RNI3L2D1_Z[0]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[0]), .FCI(GND), .S(early_val_RNIT7HB3_S[0]), .Y(
        early_val_RNIT7HB3_Y[0]), .FCO(tapcnt_final_13_m1_cry_0));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNIEOFU2[5]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[5]), .D(GND), .FCI(
        timeout_cnt_cry[4]), .S(timeout_cnt_s[5]), .Y(
        timeout_cnt_RNIEOFU2_Y[5]), .FCO(timeout_cnt_cry[5]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_153 (.A(late_flags_Z[19]), 
        .B(late_flags_Z[18]), .C(late_flags_Z[17]), .D(
        late_flags_Z[16]), .Y(calc_done25_153_Z));
    SLE \early_flags[40]  (.D(early_flags_7_fast_Z[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[40]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_180 (.A(early_flags_Z[39]), 
        .B(early_flags_Z[38]), .C(early_flags_Z[37]), .D(
        early_flags_Z[36]), .Y(calc_done25_180_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[108]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[108]), .C(
        un10_early_flags[108]), .Y(late_flags_7_fast_Z[108]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_9_1 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[9]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[31]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[31]), .C(
        un10_early_flags[31]), .Y(early_flags_7_fast_Z[31]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[12]), 
        .D(late_flags_Z[76]), .FCI(late_flags_pmux_63_1_1_co1_6), .S(
        late_flags_pmux_63_1_1_wmux_15_S), .Y(
        late_flags_pmux_63_1_1_y0_6), .FCO(
        late_flags_pmux_63_1_1_co0_7));
    SLE \early_flags[5]  (.D(early_flags_7_fast_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[5]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_130 (.A(late_flags_Z[127]), 
        .B(late_flags_Z[126]), .C(late_flags_Z[125]), .D(
        late_flags_Z[124]), .Y(calc_done25_130_Z));
    SLE \late_flags[34]  (.D(late_flags_7_fast_Z[34]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[34]));
    SLE \late_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[2])
        );
    SLE \timeout_cnt[7]  (.D(timeout_cnt_s[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[7]));
    SLE \restart_reg[2]  (.D(restart_reg_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_reg_Z[2]));
    SLE \early_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[5]));
    SLE \no_early_no_late_val_st2[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[2]));
    SLE \tapcnt_final_upd[1]  (.D(tapcnt_final_upd_8_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[1]));
    SLE \noearly_nolate_diff_nxt[7]  (.D(noearly_nolate_diff_nxt_8[7]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_7));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[26]), 
        .D(early_flags_Z[90]), .FCI(early_flags_pmux_63_1_0_co1_1), .S(
        early_flags_pmux_63_1_0_wmux_5_S), .Y(
        early_flags_pmux_63_1_0_y0_2), .FCO(
        early_flags_pmux_63_1_0_co0_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[29]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[29]), .C(
        un10_early_flags[29]), .Y(early_flags_7_fast_Z[29]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[8]), .D(
        late_flags_Z[72]), .FCI(late_flags_pmux_63_1_1_co1_0), .S(
        late_flags_pmux_63_1_1_wmux_3_S), .Y(
        late_flags_pmux_63_1_1_y0_1), .FCO(
        late_flags_pmux_63_1_1_co0_1));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_111_1_0 (.A(
        un10_early_flags_1_Z[3]), .B(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags_1_0[15]));
    CFG3 #( .INIT(8'hCD) )  rx_BIT_ALGN_DIR_0_sqmuxa_2_i (.A(
        tapcnt_final_upd_3_sqmuxa_Z), .B(restart_trng_fg_i), .C(
        un1_bitalign_curr_state_15_3_Z), .Y(
        rx_BIT_ALGN_DIR_0_sqmuxa_2_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[89]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[89]), .C(
        un10_early_flags[89]), .Y(early_flags_7_fast_Z[89]));
    SLE \early_flags[64]  (.D(early_flags_7_fast_Z[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[64]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[22]), 
        .D(early_flags_Z[86]), .FCI(early_flags_pmux_63_1_0_co1_5), .S(
        early_flags_pmux_63_1_0_wmux_13_S), .Y(
        early_flags_pmux_63_1_0_y0_5), .FCO(
        early_flags_pmux_63_1_0_co0_6));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_5 (.A(late_val_Z[5])
        , .B(early_val_Z[5]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_4_Z), .S(tapcnt_final27_cry_5_S), .Y(
        tapcnt_final27_cry_5_Y), .FCO(tapcnt_final27_cry_5_Z));
    CFG2 #( .INIT(4'h4) )  bitalign_curr_state159_2 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state159_2_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_13_1 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[5]));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[2]  (.A(
        tapcnt_final_13_Z[3]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[2]), .Y(tapcnt_final_13_1_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[63]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[63]), .C(
        un10_early_flags[63]), .Y(late_flags_7_fast_Z[63]));
    CFG2 #( .INIT(4'hE) )  un1_restart_trng_fg_10_1 (.A(
        bitalign_curr_state_1_sqmuxa_4_Z), .B(restart_trng_fg_i), .Y(
        un1_restart_trng_fg_10_sn_1));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[3]  (.A(
        tapcnt_final_13_Z[4]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[3]), .Y(tapcnt_final_13_1_Z[3]));
    SLE \early_flags[36]  (.D(early_flags_7_fast_Z[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[36]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[114]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[114]), .C(
        un10_early_flags[114]), .Y(late_flags_7_fast_Z[114]));
    SLE \late_flags[110]  (.D(late_flags_7_fast_Z[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[110]));
    SLE \early_flags[37]  (.D(early_flags_7_fast_Z[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[37]));
    SLE \early_flags[105]  (.D(early_flags_7_fast_Z[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[105]));
    SLE \early_flags[118]  (.D(early_flags_7_fast_Z[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[118]));
    CFG3 #( .INIT(8'hE4) )  \early_flags_RNO[49]  (.A(N_208), .B(
        EYE_MONITOR_EARLY_net_0_0), .C(early_flags_Z[49]), .Y(
        early_flags_RNO_Z[49]));
    CFG2 #( .INIT(4'hE) )  un1_restart_trng_fg_5 (.A(
        un1_tap_cnt_0_sqmuxa_6_0), .B(restart_trng_fg_i), .Y(
        un1_restart_trng_fg_5_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_12 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[12]));
    SLE \early_flags[120]  (.D(early_flags_7_fast_Z[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[120]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[69]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[69]), .C(
        un10_early_flags[69]), .Y(early_flags_7_fast_Z[69]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_12 (.A(
        late_flags_pmux_63_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[38]), .D(late_flags_Z[102]), .FCI(
        late_flags_pmux_63_1_0_co0_5), .S(
        late_flags_pmux_63_1_0_wmux_12_S), .Y(
        late_flags_pmux_63_1_0_y1_0), .FCO(
        late_flags_pmux_63_1_0_co1_5));
    SLE \early_flags[31]  (.D(early_flags_7_fast_Z[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[31]));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_46_3 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_3_Z[46]));
    SLE \early_flags[15]  (.D(early_flags_7_fast_Z[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[15]));
    SLE \early_flags[42]  (.D(early_flags_7_fast_Z[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[42]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_85 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[5]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[4]), .Y(
        un10_early_flags[85]));
    CFG4 #( .INIT(16'h7340) )  \bitalign_curr_state_34_4_0_.m40_1_1  (
        .A(bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[4]), .C(
        N_124_mux), .D(N_15), .Y(m40_1_1));
    SLE \noearly_nolate_diff_nxt[1]  (.D(noearly_nolate_diff_nxt_8[1]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_1));
    SLE \no_early_no_late_val_end2[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[5]));
    CFG2 #( .INIT(4'h2) )  un1_tapcnt_final (.A(un34), .B(
        un16_tapcnt_final_cry_7_Z), .Y(un1_tapcnt_final_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[5]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[5]), .C(
        un10_early_flags[5]), .Y(late_flags_7_fast_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[2]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[2]), .C(
        un10_early_flags[2]), .Y(late_flags_7_fast_Z[2]));
    SLE \early_flags[66]  (.D(early_flags_7_fast_Z[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[66]));
    CFG4 #( .INIT(16'hFFFE) )  restart_trng_fg (.A(
        restart_edge_reg_Z[3]), .B(restart_edge_reg_Z[2]), .C(
        restart_edge_reg_Z[1]), .D(restart_edge_reg_Z[0]), .Y(
        restart_trng_fg_i));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_14 (.A(
        early_flags_pmux_126_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[53]), .D(early_flags_Z[117]), .FCI(
        early_flags_pmux_126_1_1_co0_6), .S(
        early_flags_pmux_126_1_1_wmux_14_S), .Y(
        early_flags_pmux_126_1_1_y3_0), .FCO(
        early_flags_pmux_126_1_1_co1_6));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.m43_0_a2  (.A(
        bitalign_curr_state12_Z), .B(un1_rx_BIT_ALGN_START), .Y(
        bitalign_curr_state13));
    SLE \early_flags[67]  (.D(early_flags_7_fast_Z[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[67]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_2 (.A(
        early_flags_pmux_63_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[48]), .D(early_flags_Z[112]), .FCI(
        early_flags_pmux_63_1_1_co0_0), .S(
        early_flags_pmux_63_1_1_wmux_2_S), .Y(
        early_flags_pmux_63_1_1_y3), .FCO(
        early_flags_pmux_63_1_1_co1_0));
    SLE \early_flags[74]  (.D(early_flags_7_fast_Z[74]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[74]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[92]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[92]), .C(
        un10_early_flags[92]), .Y(late_flags_7_fast_Z[92]));
    CFG2 #( .INIT(4'h8) )  \bitalign_curr_state_34_4_0_.m106_1  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[3]), .Y(
        i22_mux_1));
    SLE \early_flags[119]  (.D(early_flags_7_fast_Z[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[119]));
    CFG4 #( .INIT(16'hFFEC) )  bitalign_curr_state163_RNIM5SH (.A(
        bitalign_curr_state163_Z), .B(emflag_cnt_0_sqmuxa), .C(
        bit_align_dly_done_Z), .D(restart_trng_fg_i), .Y(
        emflag_cntlde_1));
    SLE \early_flags[61]  (.D(early_flags_7_fast_Z[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[61]));
    SLE \timeout_cnt[4]  (.D(timeout_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[84]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[84]), .C(
        un10_early_flags[84]), .Y(late_flags_7_fast_Z[84]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[122]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[122]), .C(
        un10_early_flags[122]), .Y(early_flags_7_fast_Z[122]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_32_1_0_a2 (.A(tap_cnt_Z[5])
        , .B(tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[32]));
    SLE \wait_cnt[2]  (.D(wait_cnt_4_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(wait_cnt_Z[2]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_4_0 (
        .A(emflag_cnt_Z[4]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[4]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_3), .S(
        noearly_nolate_diff_start_7[4]), .Y(
        noearly_nolate_diff_start_7_cry_4_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_4));
    CFG4 #( .INIT(16'h53FF) )  \bitalign_curr_state_34_4_0_.m64_1_1  (
        .A(bitalign_curr_state41_Z), .B(N_60_0), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        m64_1_1));
    CFG1 #( .INIT(2'h1) )  un1_restart_trng_fg_5_RNIIB4C (.A(
        un1_restart_trng_fg_5_Z), .Y(N_19_i));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_126 (.A(tap_cnt_Z[0]), 
        .B(un10_early_flags_1_Z[6]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[126]));
    SLE \late_flags[82]  (.D(late_flags_7_fast_Z[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[82]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_59 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_2_Z[35]), .Y(
        un10_early_flags[59]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_35_2 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[35]));
    CFG3 #( .INIT(8'hEC) )  calc_done_0_sqmuxa_RNIFT9H (.A(
        calc_done_0_sqmuxa_Z), .B(restart_trng_fg_i), .C(
        bitalign_curr_state154_Z), .Y(timeout_cntlde_0));
    SLE \noearly_nolate_diff_nxt[0]  (.D(noearly_nolate_diff_nxt_8[0]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_0));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[113]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[113]), .C(
        un10_early_flags[113]), .Y(late_flags_7_fast_Z[113]));
    SLE \late_flags[102]  (.D(late_flags_7_fast_Z[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[102]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_87_3 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_3_Z[87]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_159 (.A(late_flags_Z[11]), 
        .B(late_flags_Z[10]), .C(late_flags_Z[9]), .D(late_flags_Z[8]), 
        .Y(calc_done25_159_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[106]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[106]), .C(
        un10_early_flags[106]), .Y(late_flags_7_fast_Z[106]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[97]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[97]), .C(
        un10_early_flags[97]), .Y(early_flags_7_fast_Z[97]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[14]), 
        .D(early_flags_Z[78]), .FCI(early_flags_pmux_63_1_0_co1_6), .S(
        early_flags_pmux_63_1_0_wmux_15_S), .Y(
        early_flags_pmux_63_1_0_y0_6), .FCO(
        early_flags_pmux_63_1_0_co0_7));
    CFG3 #( .INIT(8'h02) )  bit_align_done_2_sqmuxa (.A(
        bit_align_dly_done_0_sqmuxa_Z), .B(sig_re_train_Z), .C(
        restart_trng_fg_i), .Y(bit_align_done_2_sqmuxa_Z));
    CFG4 #( .INIT(16'h00E0) )  sig_re_train (.A(
        EYE_MONITOR_LATE_net_0_0), .B(EYE_MONITOR_EARLY_net_0_0), .C(
        un1_sig_re_train_Z), .D(BIT_ALGN_ERR_0_c), .Y(sig_re_train_Z));
    SLE \late_flags[12]  (.D(late_flags_7_fast_Z[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[12]));
    SLE \early_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[3]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_69 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[64]), .C(
        un10_early_flags_2_Z[69]), .Y(un10_early_flags[69]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_14 (.A(
        early_flags_pmux_126_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[55]), .D(early_flags_Z[119]), .FCI(
        early_flags_pmux_126_1_0_co0_6), .S(
        early_flags_pmux_126_1_0_wmux_14_S), .Y(
        early_flags_pmux_126_1_0_y3_0), .FCO(
        early_flags_pmux_126_1_0_co1_6));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_117 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_1_Z[48]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_2_Z[69]), .Y(
        un10_early_flags[117]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[56]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[56]), .C(
        un10_early_flags[56]), .Y(early_flags_7_fast_Z[56]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[72]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[72]), .C(
        un10_early_flags[72]), .Y(early_flags_7_fast_Z[72]));
    SLE \early_flags[76]  (.D(early_flags_7_fast_Z[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[76]));
    CFG4 #( .INIT(16'h0FEE) )  \bitalign_curr_state_34_4_0_.m82_1_0  (
        .A(BIT_ALGN_ERR_0_c), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .C(
        N_63), .D(bitalign_curr_state_Z[1]), .Y(m82_1_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[18]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[18]), .C(
        un10_early_flags[18]), .Y(early_flags_7_fast_Z[18]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_97 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_2_Z[69]), .D(
        un10_early_flags_2_0[96]), .Y(un10_early_flags[97]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_34 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_2_0[32]), .Y(un10_early_flags[34]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[10]), 
        .D(early_flags_Z[74]), .FCI(early_flags_pmux_63_1_0_co1_0), .S(
        early_flags_pmux_63_1_0_wmux_3_S), .Y(
        early_flags_pmux_63_1_0_y0_1), .FCO(
        early_flags_pmux_63_1_0_co0_1));
    SLE \early_flags[77]  (.D(early_flags_7_fast_Z[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[77]));
    SLE \no_early_no_late_val_end1[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[4]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_248 (.A(calc_done25_227_Z), 
        .B(calc_done25_226_Z), .C(calc_done25_225_Z), .D(
        calc_done25_224_Z), .Y(calc_done25_248_Z));
    CFG4 #( .INIT(16'h8000) )  calc_done25_229 (.A(calc_done25_151_Z), 
        .B(calc_done25_150_Z), .C(calc_done25_149_Z), .D(
        calc_done25_148_Z), .Y(calc_done25_229_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_88 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_1_Z[64]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[88]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_14 (.A(
        early_flags_pmux_63_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[54]), .D(early_flags_Z[118]), .FCI(
        early_flags_pmux_63_1_0_co0_6), .S(
        early_flags_pmux_63_1_0_wmux_14_S), .Y(
        early_flags_pmux_63_1_0_y3_0), .FCO(
        early_flags_pmux_63_1_0_co1_6));
    SLE \early_flags[111]  (.D(early_flags_7_fast_Z[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[111]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_37_2_0_a2 (.A(tap_cnt_Z[5])
        , .B(tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[37]));
    SLE \late_flags[42]  (.D(late_flags_7_fast_Z[42]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[42]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[15]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[15]), .C(
        un10_early_flags[15]), .Y(early_flags_7_fast_Z[15]));
    SLE \early_flags[71]  (.D(early_flags_7_fast_Z[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[71]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[69]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[69]), .C(
        un10_early_flags[69]), .Y(late_flags_7_fast_Z[69]));
    CFG4 #( .INIT(16'hFFFE) )  rx_BIT_ALGN_LOAD_0_sqmuxa_1_i (.A(
        restart_trng_fg_i), .B(rx_BIT_ALGN_LOAD_0_sqmuxa_Z), .C(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .D(
        un1_tap_cnt_0_sqmuxa_6_0), .Y(rx_BIT_ALGN_LOAD_0_sqmuxa_1_i_Z));
    SLE \bitalign_curr_state[4]  (.D(bitalign_curr_state_34[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[4]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_19 (.A(
        early_flags_pmux_126_1_0_y7_0), .B(
        early_flags_pmux_126_1_0_y5_0), .C(emflag_cnt_Z[4]), .D(
        emflag_cnt_Z[3]), .FCI(early_flags_pmux_126_1_0_co1_8), .S(
        early_flags_pmux_126_1_0_wmux_19_S), .Y(
        early_flags_pmux_126_1_0_y0_8), .FCO(
        early_flags_pmux_126_1_0_co0_9));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[113]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[113]), .C(
        un10_early_flags[113]), .Y(early_flags_7_fast_Z[113]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_19 (.A(
        late_flags_pmux_126_1_0_y7_0), .B(late_flags_pmux_126_1_0_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co1_8), .S(
        late_flags_pmux_126_1_0_wmux_19_S), .Y(
        late_flags_pmux_126_1_0_y0_8), .FCO(
        late_flags_pmux_126_1_0_co0_9));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_119 (.A(
        un10_early_flags_1_Z[20]), .B(tap_cnt_Z[3]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[96]), .Y(
        un10_early_flags[119]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_7 (.A(
        late_flags_pmux_126_1_0_0_y7), .B(late_flags_pmux_126_1_0_0_y5)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co1_2), .S(
        late_flags_pmux_126_1_0_wmux_7_S), .Y(
        late_flags_pmux_126_1_0_y0_3), .FCO(
        late_flags_pmux_126_1_0_co0_3));
    CFG3 #( .INIT(8'h40) )  \bitalign_curr_state_34_4_0_.m107  (.A(
        early_flags_dec[127]), .B(bitalign_curr_state89_Z), .C(
        bitalign_curr_state_Z[0]), .Y(N_108));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_24 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_2_0[24]), .C(
        un10_early_flags_1_Z[0]), .Y(un10_early_flags[24]));
    SLE \early_flags[113]  (.D(early_flags_7_fast_Z[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[113]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_2_0 (
        .A(emflag_cnt_Z[2]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[2]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_1), .S(
        noearly_nolate_diff_start_7[2]), .Y(
        noearly_nolate_diff_start_7_cry_2_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[46]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[46]), .C(
        un10_early_flags[46]), .Y(early_flags_7_fast_Z[46]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_15 (.A(
        un10_early_flags_2_0[0]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[15]));
    CFG4 #( .INIT(16'h0080) )  \bitalign_curr_state_34_4_0_.m85_2  (.A(
        bitalign_curr_state_Z[2]), .B(N_83), .C(
        bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[4]), .Y(
        m85_1));
    CFG4 #( .INIT(16'h2232) )  \bitalign_curr_state_34_4_0_.m91_1  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        un1_retrain_adj_tap_i), .D(N_69), .Y(m91_1_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[121]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[121]), .C(
        un10_early_flags[121]), .Y(early_flags_7_fast_Z[121]));
    SLE \timeout_cnt[3]  (.D(timeout_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[3]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_237 (.A(calc_done25_183_Z), 
        .B(calc_done25_182_Z), .C(calc_done25_181_Z), .D(
        calc_done25_180_Z), .Y(calc_done25_237_Z));
    CFG4 #( .INIT(16'h8000) )  calc_done25_238 (.A(calc_done25_187_Z), 
        .B(calc_done25_186_Z), .C(calc_done25_185_Z), .D(
        calc_done25_184_Z), .Y(calc_done25_238_Z));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_18 (.A(
        early_flags_pmux_63_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[62]), .D(early_flags_Z[126]), .FCI(
        early_flags_pmux_63_1_0_co0_8), .S(
        early_flags_pmux_63_1_0_wmux_18_S), .Y(
        early_flags_pmux_63_1_0_y7_0), .FCO(
        early_flags_pmux_63_1_0_co1_8));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[0]  (.A(
        un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_Y[0]), .B(N_63_0), .Y(
        N_32_i));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_107 (.A(
        un10_early_flags_1_Z[40]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_2_Z[67]), .Y(
        un10_early_flags[107]));
    SLE \timeout_cnt[1]  (.D(timeout_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[1]));
    SLE \early_flags[38]  (.D(early_flags_7_fast_Z[38]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[38]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_96 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_1_Z[96]), .C(
        un10_early_flags_2_0[96]), .Y(un10_early_flags[96]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_173 (.A(early_flags_Z[67]), 
        .B(early_flags_Z[66]), .C(early_flags_Z[65]), .D(
        early_flags_Z[64]), .Y(calc_done25_173_Z));
    SLE \late_flags[113]  (.D(late_flags_7_fast_Z[113]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[113]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[1]), .D(
        late_flags_Z[65]), .FCI(VCC), .S(
        late_flags_pmux_126_1_1_wmux_S), .Y(late_flags_pmux_126_1_1_y0)
        , .FCO(late_flags_pmux_126_1_1_co0));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[31]), 
        .D(early_flags_Z[95]), .FCI(early_flags_pmux_126_1_0_co1_7), 
        .S(early_flags_pmux_126_1_0_wmux_17_S), .Y(
        early_flags_pmux_126_1_0_y0_7), .FCO(
        early_flags_pmux_126_1_0_co0_8));
    SLE \retrain_reg[0]  (.D(sig_re_train_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(retrain_reg_Z[0]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[3]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[3]), .D(GND), .FCI(
        emflag_cnt_cry_Z[2]), .S(emflag_cnt_s[3]), .Y(
        emflag_cnt_cry_Y_0[3]), .FCO(emflag_cnt_cry_Z[3]));
    CFG4 #( .INIT(16'h0400) )  bitalign_curr_state154_3 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[2]), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state154_3_Z));
    SLE \restart_edge_reg[2]  (.D(restart_edge_reg_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[2]));
    CFG4 #( .INIT(16'h8000) )  reset_dly_fg4_6 (.A(rst_cnt_Z[5]), .B(
        rst_cnt_Z[4]), .C(rst_cnt_Z[3]), .D(rst_cnt_Z[2]), .Y(
        reset_dly_fg4_6_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[21]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[21]), .C(
        un10_early_flags[21]), .Y(early_flags_7_fast_Z[21]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_167 (.A(early_flags_Z[107]), 
        .B(early_flags_Z[106]), .C(early_flags_Z[105]), .D(
        early_flags_Z[104]), .Y(calc_done25_167_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_40_1 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_1_Z[40]));
    SLE \early_flags[29]  (.D(early_flags_7_fast_Z[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[29]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[81]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[81]), .C(
        un10_early_flags[81]), .Y(early_flags_7_fast_Z[81]));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIJGIR[1]  (.A(
        late_val_Z[1]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[1]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIJGIR_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[99]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[99]), .C(
        un10_early_flags[99]), .Y(early_flags_7_fast_Z[99]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[66]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[66]), .C(
        un10_early_flags[66]), .Y(late_flags_7_fast_Z[66]));
    CFG2 #( .INIT(4'h2) )  Restart_trng_edge_det (.A(restart_reg_Z[1]), 
        .B(restart_reg_Z[2]), .Y(Restart_trng_edge_det_Z));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_81 (.A(N_1498), .B(
        tap_cnt_Z[5]), .C(un10_early_flags_2_Z[69]), .D(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[81]));
    CFG4 #( .INIT(16'h00AC) )  \bitalign_curr_state_34_4_0_.m41  (.A(
        N_40), .B(m40_1_1), .C(bitalign_curr_state_Z[3]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[0]));
    CFG2 #( .INIT(4'h4) )  rx_BIT_ALGN_CLR_FLGS (.A(rx_trng_done_Z), 
        .B(sig_rx_BIT_ALGN_CLR_FLGS_Z), .Y(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_1_wmux_20 (.A(
        late_flags_pmux_63_1_1_y0_8), .B(late_flags_pmux_63_1_1_y3_0), 
        .C(late_flags_pmux_63_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co0_9), .S(
        late_flags_pmux_63_1_1_wmux_20_S), .Y(
        late_flags_pmux_63_1_1_y21), .FCO(late_flags_pmux_63_1_1_co1_9)
        );
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_0 (.A(
        un10_tapcnt_final_0), .B(early_late_diff_Z[0]), .C(GND), .D(
        GND), .FCI(GND), .S(un1_early_late_diff_cry_0_S), .Y(
        un1_early_late_diff_cry_0_Y), .FCO(un1_early_late_diff_cry_0_Z)
        );
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_109 (.A(
        un10_early_flags_2_Z[69]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[5]), .D(un10_early_flags_1_Z[40]), .Y(
        un10_early_flags[109]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_2 (.A(late_val_Z[2])
        , .B(early_val_Z[2]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_1_Z), .S(tapcnt_final27_cry_2_S), .Y(
        tapcnt_final27_cry_2_Y), .FCO(tapcnt_final27_cry_2_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_12_1 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[12]));
    CFG2 #( .INIT(4'h2) )  late_last_set15 (.A(early_last_set_Z), .B(
        late_last_set_Z), .Y(late_last_set15_Z));
    SLE \late_flags[111]  (.D(late_flags_7_fast_Z[111]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[111]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNO[7]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[7]), .D(GND), .FCI(
        timeout_cnt_cry[6]), .S(timeout_cnt_s[7]), .Y(
        timeout_cnt_RNO_Y[7]), .FCO(timeout_cnt_RNO_FCO[7]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_12 (.A(
        early_flags_pmux_126_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[37]), .D(early_flags_Z[101]), .FCI(
        early_flags_pmux_126_1_1_co0_5), .S(
        early_flags_pmux_126_1_1_wmux_12_S), .Y(
        early_flags_pmux_126_1_1_y1_0), .FCO(
        early_flags_pmux_126_1_1_co1_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[126]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[126]), .C(
        un10_early_flags[126]), .Y(late_flags_7_fast_Z[126]));
    CFG2 #( .INIT(4'h8) )  calc_done_4_sqmuxa_0 (.A(
        bitalign_curr_state162_Z), .B(un1_early_late_diff_valid_Z), .Y(
        calc_done_4_sqmuxa_0_Z));
    SLE \late_flags[92]  (.D(late_flags_7_fast_Z[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[92]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[61]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[61]), .C(
        un10_early_flags[61]), .Y(early_flags_7_fast_Z[61]));
    SLE \early_flags[68]  (.D(early_flags_7_fast_Z[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[68]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_11_1 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_1_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[94]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[94]), .C(
        un10_early_flags[94]), .Y(late_flags_7_fast_Z[94]));
    SLE \bitalign_curr_state[0]  (.D(bitalign_curr_state_34[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[0]));
    CFG2 #( .INIT(4'h8) )  bitalign_curr_state152_1 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[1]), .Y(
        bitalign_curr_state152_1_Z));
    CFG2 #( .INIT(4'h2) )  rx_BIT_ALGN_START (.A(bit_align_start_Z), 
        .B(BIT_ALGN_ERR_0_c), .Y(BIT_ALGN_START_1_c));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[51]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[51]), .C(
        un10_early_flags[51]), .Y(late_flags_7_fast_Z[51]));
    CFG3 #( .INIT(8'h40) )  bitalign_curr_state159 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state159_2_Z), .C(
        bitalign_curr_state155_1_Z), .Y(bitalign_curr_state159_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[0]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[0]), .C(
        un10_early_flags[0]), .Y(early_flags_7_fast_Z[0]));
    CFG4 #( .INIT(16'h331B) )  \bitalign_curr_state_34_4_0_.m23  (.A(
        N_117_mux_1), .B(bitalign_curr_state_Z[1]), .C(m23_1_2), .D(
        early_flags_dec[127]), .Y(N_124_mux));
    CFG3 #( .INIT(8'h40) )  un10_early_flags_18 (.A(N_1499), .B(
        un10_early_flags_2_Z[10]), .C(un10_early_flags_2_0[16]), .Y(
        un10_early_flags[18]));
    CFG4 #( .INIT(16'hEFEE) )  un1_bitalign_curr_state_0_sqmuxa_9_1 (
        .A(early_flags_0_sqmuxa_Z), .B(
        bitalign_curr_state_0_sqmuxa_8_Z), .C(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .D(bitalign_curr_state154_Z), 
        .Y(un1_bitalign_curr_state_0_sqmuxa_9_1_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_165 (.A(early_flags_Z[99]), 
        .B(early_flags_Z[98]), .C(early_flags_Z[97]), .D(
        early_flags_Z[96]), .Y(calc_done25_165_Z));
    CFG4 #( .INIT(16'hFFFE) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i (
        .A(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .B(
        un1_bitalign_curr_state_1_sqmuxa_6_i_0), .C(restart_trng_fg_i), 
        .D(un1_rx_BIT_ALGN_LOAD_0_sqmuxa_i_0), .Y(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i_Z));
    SLE \late_flags[56]  (.D(late_flags_7_fast_Z[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[56]));
    SLE \early_flags[102]  (.D(early_flags_7_fast_Z[102]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[102]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIP2921[0]  (.A(
        no_early_no_late_val_st1_Z[0]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[0]), .Y(
        un1_no_early_no_late_val_st1_1_1[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_2 (.A(
        late_flags_pmux_63_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[48]), .D(late_flags_Z[112]), .FCI(
        late_flags_pmux_63_1_1_co0_0), .S(
        late_flags_pmux_63_1_1_wmux_2_S), .Y(late_flags_pmux_63_1_1_y3)
        , .FCO(late_flags_pmux_63_1_1_co1_0));
    SLE \late_flags[20]  (.D(late_flags_7_fast_Z[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[20]));
    CFG3 #( .INIT(8'h20) )  early_last_set_1_sqmuxa_1_3 (.A(N_20), .B(
        late_last_set15_Z), .C(bitalign_curr_state161_Z), .Y(
        early_last_set_1_sqmuxa_1_3_Z));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_1_wmux_20 (.A(
        early_flags_pmux_126_1_1_y0_8), .B(
        early_flags_pmux_126_1_1_y3_0), .C(
        early_flags_pmux_126_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_1_co0_9), .S(
        early_flags_pmux_126_1_1_wmux_20_S), .Y(
        early_flags_pmux_126_1_1_y21), .FCO(
        early_flags_pmux_126_1_1_co1_9));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_8 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[3]), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[8]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[127]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[127]), .C(
        un10_early_flags[127]), .Y(early_flags_7_fast_Z[127]));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_80 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[0]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[0]), .Y(
        un10_early_flags[80]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_1_0 (.A(
        emflag_cnt_Z[1]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[1]), .D(GND), .FCI(early_late_diff_8_cry_0), .S(
        early_late_diff_8[1]), .Y(early_late_diff_8_cry_1_0_Y), .FCO(
        early_late_diff_8_cry_1));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_2 (.A(
        un16_tapcnt_final_2), .B(un10_tapcnt_final_2), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_1_Z), .S(
        un16_tapcnt_final_cry_2_S), .Y(un16_tapcnt_final_cry_2_Y), 
        .FCO(un16_tapcnt_final_cry_2_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_9 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_126_1_0_co1_3), .S(
        early_flags_pmux_126_1_0_wmux_9_S), .Y(
        early_flags_pmux_126_1_0_wmux_9_Y), .FCO(
        early_flags_pmux_126_1_0_co0_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[77]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[77]), .C(
        un10_early_flags[77]), .Y(early_flags_7_fast_Z[77]));
    CFG4 #( .INIT(16'h00CE) )  \bitalign_curr_state_34_4_0_.m86  (.A(
        m86_1), .B(m85_1), .C(bitalign_curr_state_Z[3]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[2]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_2 (.A(
        late_flags_pmux_126_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[49]), .D(late_flags_Z[113]), .FCI(
        late_flags_pmux_126_1_1_co0_0), .S(
        late_flags_pmux_126_1_1_wmux_2_S), .Y(
        late_flags_pmux_126_1_1_y3), .FCO(
        late_flags_pmux_126_1_1_co1_0));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[109]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[109]), .C(
        un10_early_flags[109]), .Y(late_flags_7_fast_Z[109]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[13]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[13]), .C(
        un10_early_flags[13]), .Y(early_flags_7_fast_Z[13]));
    CFG4 #( .INIT(16'h08FF) )  un1_early_flags_pmux_1_RNI26QC (.A(
        late_last_set15_Z), .B(bitalign_curr_state161_Z), .C(
        un1_early_flags_pmux_1_Z), .D(early_late_diff_0_sqmuxa_1_0_Z), 
        .Y(no_early_no_late_val_end2_0_sqmuxa_i));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_37 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[32]), .C(
        un10_early_flags_2_Z[37]), .Y(un10_early_flags[37]));
    SLE \tap_cnt[6]  (.D(N_1496_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tap_cnt_Z[6]));
    CFG2 #( .INIT(4'hE) )  rx_BIT_ALGN_DONE (.A(bit_align_done_Z), .B(
        BIT_ALGN_ERR_0_c), .Y(BIT_ALGN_DONE_c));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_10 (.A(
        late_flags_pmux_126_1_0_0_y21), .B(
        late_flags_pmux_126_1_0_0_y9), .C(emflag_cnt_Z[2]), .D(VCC), 
        .FCI(late_flags_pmux_126_1_0_co0_4), .S(
        late_flags_pmux_126_1_0_wmux_10_S), .Y(
        late_flags_pmux_126_1_0_wmux_10_Y), .FCO(
        late_flags_pmux_126_1_0_co1_4));
    SLE \early_flags[78]  (.D(early_flags_7_fast_Z[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[78]));
    CFG3 #( .INIT(8'h08) )  tapcnt_final_upd_2_sqmuxa_0_a2 (.A(
        mv_up_fg_Z), .B(N_100), .C(mv_dn_fg_Z), .Y(
        tapcnt_final_upd_2_sqmuxa));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_0 (.A(
        early_flags_pmux_63_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[34]), .D(early_flags_Z[98]), .FCI(
        early_flags_pmux_63_1_0_0_co0), .S(
        early_flags_pmux_63_1_0_wmux_0_S), .Y(
        early_flags_pmux_63_1_0_0_y1), .FCO(
        early_flags_pmux_63_1_0_0_co1));
    CFG4 #( .INIT(16'h3AFA) )  \bitalign_curr_state_34_4_0_.m67_1  (.A(
        N_51), .B(N_119_mux), .C(bitalign_curr_state_Z[4]), .D(m55_0), 
        .Y(m67_1));
    SLE \late_flags[70]  (.D(late_flags_7_fast_Z[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[70]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_48_2_0 (.A(
        un10_early_flags_2_Z[0]), .B(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[48]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_3_0 (.A(
        emflag_cnt_Z[3]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[3]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_2), .S(
        noearly_nolate_diff_nxt_8[3]), .Y(
        noearly_nolate_diff_nxt_8_cry_3_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_3));
    SLE \noearly_nolate_diff_start[0]  (.D(
        noearly_nolate_diff_start_7[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_0));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_42 (.A(
        un10_early_flags_1_Z[10]), .B(un10_early_flags_1_Z[32]), .C(
        un10_early_flags_2_0[40]), .Y(un10_early_flags[42]));
    CFG3 #( .INIT(8'hFD) )  rx_BIT_ALGN_MOVE_0_sqmuxa_2_i (.A(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_1_Z), .B(
        un1_restart_trng_fg_10_sn_1), .C(tap_cnt_0_sqmuxa_1_Z), .Y(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_i_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_147 (.A(late_flags_Z[55]), 
        .B(late_flags_Z[54]), .C(late_flags_Z[53]), .D(
        late_flags_Z[52]), .Y(calc_done25_147_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[71]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[71]), .C(
        un10_early_flags[71]), .Y(late_flags_7_fast_Z[71]));
    SLE \no_early_no_late_val_end2[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[2]));
    SLE \late_flags[66]  (.D(late_flags_7_fast_Z[66]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[66]));
    CFG4 #( .INIT(16'h1101) )  \bitalign_curr_state_34_4_0_.m37_0  (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[0]), .C(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .D(BIT_ALGN_ERR_0_c), .Y(m37));
    ARI1 #( .INIT(20'h44844) )  tapcnt_final_upd_8_s_6 (.A(N_100), .B(
        tap_cnt_Z[6]), .C(N_12_i), .D(mv_up_fg_Z), .FCI(
        tapcnt_final_upd_8_cry_5), .S(tapcnt_final_upd_8[6]), .Y(
        tapcnt_final_upd_8_s_6_Y), .FCO(tapcnt_final_upd_8_s_6_FCO));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_12 (.A(
        early_flags_pmux_63_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[36]), .D(early_flags_Z[100]), .FCI(
        early_flags_pmux_63_1_1_co0_5), .S(
        early_flags_pmux_63_1_1_wmux_12_S), .Y(
        early_flags_pmux_63_1_1_y1_0), .FCO(
        early_flags_pmux_63_1_1_co1_5));
    CFG4 #( .INIT(16'h0001) )  calc_done25_179 (.A(early_flags_Z[59]), 
        .B(early_flags_Z[58]), .C(early_flags_Z[57]), .D(
        early_flags_Z[56]), .Y(calc_done25_179_Z));
    CFG3 #( .INIT(8'hEA) )  un2_noearly_nolate_diff_start_validlto2 (
        .A(un10_tapcnt_final_2), .B(un10_tapcnt_final_1), .C(
        un10_tapcnt_final_0), .Y(
        un2_noearly_nolate_diff_start_validlt3));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[4]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[4]), .C(
        un10_early_flags[4]), .Y(early_flags_7_fast_Z[4]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_251 (.A(calc_done25_239_Z), 
        .B(calc_done25_238_Z), .C(calc_done25_237_Z), .D(
        calc_done25_236_Z), .Y(calc_done25_251_Z));
    SLE \tapcnt_final[3]  (.D(tapcnt_final_13_1_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[3]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_10 (.A(
        early_flags_pmux_126_1_0_0_y21), .B(
        early_flags_pmux_126_1_0_0_y9), .C(emflag_cnt_Z[2]), .D(VCC), 
        .FCI(early_flags_pmux_126_1_0_co0_4), .S(
        early_flags_pmux_126_1_0_wmux_10_S), .Y(
        early_flags_pmux_126_1_0_wmux_10_Y), .FCO(
        early_flags_pmux_126_1_0_co1_4));
    CFG2 #( .INIT(4'h8) )  bitalign_curr_state152_3 (.A(
        bitalign_curr_state152_1_Z), .B(bitalign_curr_state148_2_Z), 
        .Y(bitalign_curr_state152_3_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_27 (.A(
        un10_early_flags_2_0[24]), .B(un10_early_flags_1_Z[24]), .C(
        un10_early_flags_1_Z[3]), .Y(un10_early_flags[27]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_11 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[11]));
    CFG4 #( .INIT(16'hFFC8) )  un1_bitalign_curr_state_0_sqmuxa_9_4 (
        .A(calc_done28_Z), .B(bitalign_curr_state162_Z), .C(
        calc_done27_Z), .D(un1_bitalign_curr_state_0_sqmuxa_9_2_Z), .Y(
        un1_bitalign_curr_state_0_sqmuxa_9_4_Z));
    SLE \bitalign_curr_state[3]  (.D(bitalign_curr_state_34[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[3]));
    SLE \tapcnt_final_upd[3]  (.D(tapcnt_final_upd_8[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[3]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_120 (.A(tap_cnt_Z[2]), 
        .B(un10_early_flags_1_Z[0]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[120]));
    SLE \late_flags[30]  (.D(late_flags_7_fast_Z[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[30]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_73 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_Z[69]), .C(
        un10_early_flags_2_0[72]), .Y(un10_early_flags[73]));
    SLE \late_flags[51]  (.D(late_flags_7_fast_Z[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[51]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[9]), 
        .D(early_flags_Z[73]), .FCI(early_flags_pmux_126_1_1_co1_0), 
        .S(early_flags_pmux_126_1_1_wmux_3_S), .Y(
        early_flags_pmux_126_1_1_y0_1), .FCO(
        early_flags_pmux_126_1_1_co0_1));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_0 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[53]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[53]), .C(
        un10_early_flags[53]), .Y(late_flags_7_fast_Z[53]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_6 (.A(
        un10_tapcnt_final_6), .B(early_late_diff_Z[6]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_5_Z), .S(
        un1_early_late_diff_cry_6_S), .Y(un1_early_late_diff_cry_6_Y), 
        .FCO(un1_early_late_diff_cry_6_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_187 (.A(early_flags_Z[27]), 
        .B(early_flags_Z[26]), .C(early_flags_Z[25]), .D(
        early_flags_Z[24]), .Y(calc_done25_187_Z));
    CFG2 #( .INIT(4'h1) )  rx_trng_done1_2_sqmuxa_0_398_i_a5 (.A(
        mv_up_fg_Z), .B(mv_dn_fg_Z), .Y(N_1416));
    CFG4 #( .INIT(16'h2000) )  tapcnt_final_3_sqmuxa (.A(
        bitalign_curr_state162_Z), .B(un1_calc_done25_5_Z), .C(
        tapcnt_final27), .D(un1_early_late_diff_valid_Z), .Y(
        tapcnt_final_3_sqmuxa_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_6 (.A(
        late_flags_pmux_126_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[59]), .D(late_flags_Z[123]), .FCI(
        late_flags_pmux_126_1_0_co0_2), .S(
        late_flags_pmux_126_1_0_wmux_6_S), .Y(
        late_flags_pmux_126_1_0_0_y7), .FCO(
        late_flags_pmux_126_1_0_co1_2));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_36 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_2_0[32]), .C(
        un10_early_flags_1_Z[36]), .Y(un10_early_flags[36]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[32]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[32]), .C(
        un10_early_flags[32]), .Y(late_flags_7_fast_Z[32]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[0]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[0]), .D(GND), .FCI(
        emflag_cnt_cry_cy), .S(emflag_cnt_s[0]), .Y(
        emflag_cnt_cry_Y_0[0]), .FCO(emflag_cnt_cry_Z[0]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_137 (.A(late_flags_Z[83]), 
        .B(late_flags_Z[82]), .C(late_flags_Z[81]), .D(
        late_flags_Z[80]), .Y(calc_done25_137_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_150 (.A(late_flags_Z[47]), 
        .B(late_flags_Z[46]), .C(late_flags_Z[45]), .D(
        late_flags_Z[44]), .Y(calc_done25_150_Z));
    CFG2 #( .INIT(4'h8) )  \tapcnt_final_13_1[6]  (.A(
        tapcnt_final_13_Z[6]), .B(un1_tapcnt_final_0_sqmuxa_Z), .Y(
        tapcnt_final_13_1_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[20]), 
        .D(late_flags_Z[84]), .FCI(late_flags_pmux_63_1_1_co1_5), .S(
        late_flags_pmux_63_1_1_wmux_13_S), .Y(
        late_flags_pmux_63_1_1_y0_5), .FCO(
        late_flags_pmux_63_1_1_co0_6));
    SLE \early_flags[115]  (.D(early_flags_7_fast_Z[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[115]));
    SLE \late_flags[117]  (.D(late_flags_7_fast_Z[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[117]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[103]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[103]), .C(
        un10_early_flags[103]), .Y(early_flags_7_fast_Z[103]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[15]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[15]), .C(
        un10_early_flags[15]), .Y(late_flags_7_fast_Z[15]));
    SLE \tapcnt_final[4]  (.D(tapcnt_final_13_1_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[22]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[22]), .C(
        un10_early_flags[22]), .Y(late_flags_7_fast_Z[22]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[19]), 
        .D(early_flags_Z[83]), .FCI(early_flags_pmux_126_1_0_0_co1), 
        .S(early_flags_pmux_126_1_0_wmux_1_S), .Y(
        early_flags_pmux_126_1_0_y0_0), .FCO(
        early_flags_pmux_126_1_0_co0_0));
    SLE \no_early_no_late_val_st1[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[1]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_145 (.A(late_flags_Z[59]), 
        .B(late_flags_Z[58]), .C(late_flags_Z[57]), .D(
        late_flags_Z[56]), .Y(calc_done25_145_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_20_1 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[20]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_116 (.A(tap_cnt_Z[3]), 
        .B(un10_early_flags_1_Z[20]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[116]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[79]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[79]), .C(
        un10_early_flags[79]), .Y(early_flags_7_fast_Z[79]));
    CFG2 #( .INIT(4'h2) )  early_flags_1_sqmuxa (.A(
        bitalign_curr_state153_Z), .B(BIT_ALGN_OOR_c), .Y(
        early_flags_1_sqmuxa_Z));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_1 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[0]), .D(
        un10_early_flags_2_Z[0]), .Y(un10_early_flags[1]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_7 (.A(
        late_flags_pmux_63_1_1_y7), .B(late_flags_pmux_63_1_1_y5), .C(
        emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co1_2), .S(
        late_flags_pmux_63_1_1_wmux_7_S), .Y(
        late_flags_pmux_63_1_1_y0_3), .FCO(
        late_flags_pmux_63_1_1_co0_3));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_26 (.A(
        un10_early_flags_1_Z[10]), .B(un10_early_flags_2_0[24]), .C(
        un10_early_flags_1_Z[16]), .Y(un10_early_flags[26]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_10 (.A(
        un10_early_flags_1_Z[10]), .B(un10_early_flags_2_Z[10]), .C(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[10]));
    SLE \late_flags[61]  (.D(late_flags_7_fast_Z[61]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[61]));
    SLE \early_flags[14]  (.D(early_flags_7_fast_Z[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[14]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNI3D921[5]  (.A(
        no_early_no_late_val_st1_Z[5]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[5]), .Y(
        un1_no_early_no_late_val_st1_1_1[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[91]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[91]), .C(
        un10_early_flags[91]), .Y(early_flags_7_fast_Z[91]));
    CFG3 #( .INIT(8'hB1) )  \bitalign_curr_state_34_4_0_.m14  (.A(
        bitalign_curr_state_Z[2]), .B(N_8), .C(N_14), .Y(N_15));
    CFG4 #( .INIT(16'h0001) )  calc_done25_185 (.A(early_flags_Z[19]), 
        .B(early_flags_Z[18]), .C(early_flags_Z[17]), .D(
        early_flags_Z[16]), .Y(calc_done25_185_Z));
    CFG4 #( .INIT(16'h0CAE) )  un1_bitalign_curr_state148_9_0 (.A(
        bitalign_curr_state154_Z), .B(bitalign_curr_state164_Z), .C(
        bitalign_curr_state41_Z), .D(calc_done_0_sqmuxa_Z), .Y(
        un1_bitalign_curr_state148_9_0_Z));
    ARI1 #( .INIT(20'h4AA00) )  rst_cnt_s_715 (.A(VCC), .B(
        rst_cnt_Z[0]), .C(GND), .D(GND), .FCI(VCC), .S(rst_cnt_s_715_S)
        , .Y(rst_cnt_s_715_Y), .FCO(rst_cnt_s_715_FCO));
    SLE \no_early_no_late_val_st2[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[110]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[110]), .C(
        un10_early_flags[110]), .Y(late_flags_7_fast_Z[110]));
    SLE \rst_cnt[3]  (.D(rst_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[73]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[73]), .C(
        un10_early_flags[73]), .Y(late_flags_7_fast_Z[73]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[42]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[42]), .C(
        un10_early_flags[42]), .Y(late_flags_7_fast_Z[42]));
    SLE \late_flags[25]  (.D(late_flags_7_fast_Z[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[25]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[110]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[110]), .C(
        un10_early_flags[110]), .Y(early_flags_7_fast_Z[110]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_135 (.A(late_flags_Z[107]), 
        .B(late_flags_Z[106]), .C(late_flags_Z[105]), .D(
        late_flags_Z[104]), .Y(calc_done25_135_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_2 (.A(
        un16_tapcnt_final_2), .B(early_late_diff_Z[2]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_1_Z), .S(
        un1_early_late_diff_1_cry_2_S), .Y(
        un1_early_late_diff_1_cry_2_Y), .FCO(
        un1_early_late_diff_1_cry_2_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[10]), 
        .D(late_flags_Z[74]), .FCI(late_flags_pmux_63_1_0_co1_0), .S(
        late_flags_pmux_63_1_0_wmux_3_S), .Y(
        late_flags_pmux_63_1_0_y0_1), .FCO(
        late_flags_pmux_63_1_0_co0_1));
    SLE \early_flags[49]  (.D(early_flags_RNO_Z[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[49]));
    CFG4 #( .INIT(16'h8000) )  rx_BIT_ALGN_ERR_4 (.A(timeout_cnt_Z[3]), 
        .B(timeout_cnt_Z[2]), .C(timeout_cnt_Z[1]), .D(
        timeout_cnt_Z[0]), .Y(rx_BIT_ALGN_ERR_4_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[7]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[7]), .C(
        un10_early_flags[7]), .Y(late_flags_7_fast_Z[7]));
    ARI1 #( .INIT(20'h574B8) )  \tapcnt_final_RNIC3R56[5]  (.A(
        tap_cnt_Z[5]), .B(un1_tap_cnt_0_sqmuxa_14_0_Z[1]), .C(N_60), 
        .D(tapcnt_final_Z[5]), .FCI(tap_cnt_17_i_m2_cry_4), .S(N_75), 
        .Y(tapcnt_final_RNIC3R56_Y[5]), .FCO(tap_cnt_17_i_m2_cry_5));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[4]  (.A(N_76), .B(N_63_0), .Y(
        N_24_i));
    SLE \noearly_nolate_diff_nxt[4]  (.D(noearly_nolate_diff_nxt_8[4]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_4));
    SLE \late_flags[106]  (.D(late_flags_7_fast_Z[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[106]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_45 (.A(
        un10_early_flags_2_0[44]), .B(un10_early_flags_1_Z[40]), .C(
        un10_early_flags_1_Z[5]), .Y(un10_early_flags[45]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_106 (.A(
        un10_early_flags_1_Z[10]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[96]), .D(un10_early_flags_2_Z[10]), .Y(
        un10_early_flags[106]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[115]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[115]), .C(
        un10_early_flags[115]), .Y(late_flags_7_fast_Z[115]));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_1_wmux_8 (.A(
        early_flags_pmux_126_1_1_y0_3), .B(early_flags_pmux_126_1_1_y3)
        , .C(early_flags_pmux_126_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_1_co0_3), .S(
        early_flags_pmux_126_1_1_wmux_8_S), .Y(
        early_flags_pmux_126_1_1_y9), .FCO(
        early_flags_pmux_126_1_1_co1_3));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_0_wmux_7 (.A(
        early_flags_pmux_126_1_0_0_y7), .B(
        early_flags_pmux_126_1_0_0_y5), .C(emflag_cnt_Z[4]), .D(
        emflag_cnt_Z[3]), .FCI(early_flags_pmux_126_1_0_co1_2), .S(
        early_flags_pmux_126_1_0_wmux_7_S), .Y(
        early_flags_pmux_126_1_0_y0_3), .FCO(
        early_flags_pmux_126_1_0_co0_3));
    SLE \early_flags[16]  (.D(early_flags_7_fast_Z[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[16]));
    SLE \tapcnt_final[2]  (.D(tapcnt_final_13_1_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[2]));
    SLE \late_flags[87]  (.D(late_flags_7_fast_Z[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[87]));
    SLE \early_flags[17]  (.D(early_flags_7_fast_Z[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[17]));
    CFG2 #( .INIT(4'hE) )  \tap_cnt_17_i_o2[6]  (.A(
        un1_bitalign_curr_state_1_sqmuxa_2_i_0), .B(restart_trng_fg_i), 
        .Y(N_63_0));
    CFG3 #( .INIT(8'h80) )  calc_done_0_sqmuxa (.A(calc_done_Z), .B(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .C(rx_err_Z), .Y(
        calc_done_0_sqmuxa_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[107]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[107]), .C(
        un10_early_flags[107]), .Y(late_flags_7_fast_Z[107]));
    SLE \early_flags[33]  (.D(early_flags_7_fast_Z[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[33]));
    CFG4 #( .INIT(16'hECFE) )  un1_bitalign_curr_state_15_0 (.A(
        bitalign_curr_state_Z[1]), .B(un1_bitalign_curr_state_15_1_Z), 
        .C(bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state_15_0_Z));
    SLE late_last_set (.D(early_late_diff_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(late_last_set_Z));
    SLE \late_flags[75]  (.D(late_flags_7_fast_Z[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[75]));
    CFG2 #( .INIT(4'h2) )  late_cur_set_2_sqmuxa (.A(
        un1_bitalign_curr_state_2_sqmuxa_Z), .B(restart_trng_fg_i), .Y(
        late_cur_set_2_sqmuxa_Z));
    CFG2 #( .INIT(4'h8) )  rx_BIT_ALGN_MOVE_0_sqmuxa_1 (.A(
        bitalign_curr_state156_Z), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z));
    SLE \early_flags[50]  (.D(early_flags_RNO_Z[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[50]));
    CFG4 #( .INIT(16'h5504) )  \bitalign_curr_state_34_4_0_.m93  (.A(
        early_flags_dec[127]), .B(N_20), .C(late_last_set15_Z), .D(
        bitalign_curr_state_Z[0]), .Y(N_94));
    CFG2 #( .INIT(4'h1) )  
        \bitalign_curr_state148.bitalign_curr_state148_3_1  (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state163_2));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_0_wmux_20 (.A(
        early_flags_pmux_63_1_0_y0_8), .B(early_flags_pmux_63_1_0_y3_0)
        , .C(early_flags_pmux_63_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co0_9), .S(
        early_flags_pmux_63_1_0_wmux_20_S), .Y(
        early_flags_pmux_63_1_0_0_y21), .FCO(
        early_flags_pmux_63_1_0_co1_9));
    SLE \early_flags[11]  (.D(early_flags_7_fast_Z[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[11]));
    CFG4 #( .INIT(16'hFFC8) )  un1_bitalign_curr_state_0_sqmuxa_9_2 (
        .A(calc_done25_Z), .B(bitalign_curr_state162_Z), .C(
        calc_done26_Z), .D(un1_bitalign_curr_state_0_sqmuxa_9_1_Z), .Y(
        un1_bitalign_curr_state_0_sqmuxa_9_2_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_3 (.A(
        un16_tapcnt_final_3), .B(early_late_diff_Z[3]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_2_Z), .S(
        un1_early_late_diff_1_cry_3_S), .Y(
        un1_early_late_diff_1_cry_3_Y), .FCO(
        un1_early_late_diff_1_cry_3_Z));
    SLE \no_early_no_late_val_end1[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[1]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[24]), 
        .D(early_flags_Z[88]), .FCI(early_flags_pmux_63_1_1_co1_1), .S(
        early_flags_pmux_63_1_1_wmux_5_S), .Y(
        early_flags_pmux_63_1_1_y0_2), .FCO(
        early_flags_pmux_63_1_1_co0_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[30]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[30]), .C(
        un10_early_flags[30]), .Y(early_flags_7_fast_Z[30]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[59]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[59]), .C(
        un10_early_flags[59]), .Y(late_flags_7_fast_Z[59]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_4 (.A(
        un10_tapcnt_final_4), .B(un16_tapcnt_final_4), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_3_Z), .S(
        un10_tapcnt_final_cry_4_S), .Y(un10_tapcnt_final_cry_4_Y), 
        .FCO(un10_tapcnt_final_cry_4_Z));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_5 (.A(
        tapcnt_final_upd_Z[5]), .B(tapcnt_final_Z[5]), .C(tap_cnt_Z[5])
        , .D(N_1416), .Y(bitalign_curr_state61_5_Z));
    SLE \late_flags[17]  (.D(late_flags_7_fast_Z[17]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[17]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[17]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[17]), .C(
        un10_early_flags[17]), .Y(late_flags_7_fast_Z[17]));
    SLE \tapcnt_final[0]  (.D(tapcnt_final_13_1_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[18]), 
        .D(early_flags_Z[82]), .FCI(early_flags_pmux_63_1_0_0_co1), .S(
        early_flags_pmux_63_1_0_wmux_1_S), .Y(
        early_flags_pmux_63_1_0_y0_0), .FCO(
        early_flags_pmux_63_1_0_co0_0));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_84 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[64]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[4]), .Y(
        un10_early_flags[84]));
    SLE \late_flags[35]  (.D(late_flags_7_fast_Z[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[35]));
    SLE \early_flags[25]  (.D(early_flags_7_fast_Z[25]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[25]));
    CFG4 #( .INIT(16'h1302) )  \bitalign_curr_state_34_4_0_.m39  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[4]), .C(
        i12_mux_0), .D(N_31), .Y(N_40));
    CFG4 #( .INIT(16'hF0CA) )  \bitalign_curr_state_34_4_0_.m74_1_0  (
        .A(N_9), .B(N_11), .C(rx_err_Z), .D(bitalign_curr_state_Z[1]), 
        .Y(m74_1_0));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_1_0 (.A(
        emflag_cnt_Z[1]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[1]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_0), .S(
        noearly_nolate_diff_nxt_8[1]), .Y(
        noearly_nolate_diff_nxt_8_cry_1_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_1));
    CFG4 #( .INIT(16'h8000) )  calc_done25_249 (.A(calc_done25_231_Z), 
        .B(calc_done25_230_Z), .C(calc_done25_229_Z), .D(
        calc_done25_228_Z), .Y(calc_done25_249_Z));
    SLE \early_flags[63]  (.D(early_flags_7_fast_Z[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[63]));
    SLE \rst_cnt[6]  (.D(rst_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[6]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_118 (.A(tap_cnt_Z[3]), 
        .B(un10_early_flags_1_Z[6]), .C(un10_early_flags_1_Z[64]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[118]));
    CFG2 #( .INIT(4'h4) )  \tapcnt_final_upd_8[0]  (.A(
        mv_dn_fg_0_sqmuxa_i_o2_Z), .B(tap_cnt_Z[0]), .Y(
        tapcnt_final_upd_8_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[52]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[52]), .C(
        un10_early_flags[52]), .Y(early_flags_7_fast_Z[52]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[31]), 
        .D(late_flags_Z[95]), .FCI(late_flags_pmux_126_1_0_co1_7), .S(
        late_flags_pmux_126_1_0_wmux_17_S), .Y(
        late_flags_pmux_126_1_0_y0_7), .FCO(
        late_flags_pmux_126_1_0_co0_8));
    SLE \late_flags[47]  (.D(late_flags_7_fast_Z[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[47]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_4 (.A(
        un16_tapcnt_final_4), .B(early_late_diff_Z[4]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_3_Z), .S(
        un1_early_late_diff_1_cry_4_S), .Y(
        un1_early_late_diff_1_cry_4_Y), .FCO(
        un1_early_late_diff_1_cry_4_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_52 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[32]), .C(
        un10_early_flags_2_0[52]), .Y(un10_early_flags[52]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_10 (.A(
        late_flags_pmux_126_1_1_y21), .B(late_flags_pmux_126_1_1_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_126_1_1_co0_4), .S(
        late_flags_pmux_126_1_1_wmux_10_S), .Y(
        late_flags_pmux_126_1_1_wmux_10_Y), .FCO(
        late_flags_pmux_126_1_1_co1_4));
    SLE \emflag_cnt[4]  (.D(emflag_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[34]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[34]), .C(
        un10_early_flags[34]), .Y(late_flags_7_fast_Z[34]));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state148_5 (.A(
        bitalign_curr_state162_Z), .B(un1_bitalign_curr_state148_5_4_Z)
        , .C(bitalign_curr_state164_Z), .Y(
        un1_bitalign_curr_state148_5_Z));
    CFG3 #( .INIT(8'h80) )  calc_done25 (.A(calc_done25_248_Z), .B(
        calc_done25_253_Z), .C(calc_done25_249_Z), .Y(calc_done25_Z));
    SLE \late_flags[1]  (.D(late_flags_7_fast_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[1]));
    CFG3 #( .INIT(8'hE4) )  \early_flags_RNO[50]  (.A(N_209), .B(
        EYE_MONITOR_EARLY_net_0_0), .C(early_flags_Z[50]), .Y(
        early_flags_RNO_Z[50]));
    CFG4 #( .INIT(16'h4073) )  \bitalign_curr_state_34_4_0_.m7_1_0  (
        .A(BIT_ALGN_OOR_c), .B(bitalign_curr_state_Z[0]), .C(
        bitalign_curr_state41_Z), .D(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .Y(
        m7_1_1));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_14 (.A(
        late_flags_pmux_63_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[54]), .D(late_flags_Z[118]), .FCI(
        late_flags_pmux_63_1_0_co0_6), .S(
        late_flags_pmux_63_1_0_wmux_14_S), .Y(
        late_flags_pmux_63_1_0_y3_0), .FCO(
        late_flags_pmux_63_1_0_co1_6));
    CFG2 #( .INIT(4'hE) )  un1_sig_re_train (.A(rx_trng_done_Z), .B(
        rx_trng_done1_Z), .Y(un1_sig_re_train_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_1 (.A(
        un16_tapcnt_final_1), .B(early_late_diff_Z[1]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_0_Z), .S(
        un1_early_late_diff_1_cry_1_S), .Y(
        un1_early_late_diff_1_cry_1_Y), .FCO(
        un1_early_late_diff_1_cry_1_Z));
    SLE \early_flags[106]  (.D(early_flags_7_fast_Z[106]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[106]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[24]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[24]), .C(
        un10_early_flags[24]), .Y(late_flags_7_fast_Z[24]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_12 (.A(
        late_flags_pmux_63_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[36]), .D(late_flags_Z[100]), .FCI(
        late_flags_pmux_63_1_1_co0_5), .S(
        late_flags_pmux_63_1_1_wmux_12_S), .Y(
        late_flags_pmux_63_1_1_y1_0), .FCO(
        late_flags_pmux_63_1_1_co1_5));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIROIR[5]  (.A(
        late_val_Z[5]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[5]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIROIR_Z[5]));
    SLE \early_flags[52]  (.D(early_flags_7_fast_Z[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[52]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_48 (.A(
        un10_early_flags_1_Z[0]), .B(un10_early_flags_1_Z[48]), .C(
        un10_early_flags_2_0[48]), .Y(un10_early_flags[48]));
    CFG2 #( .INIT(4'h2) )  tap_cnt_0_sqmuxa_1_0 (.A(
        tap_cnt_0_sqmuxa_0_Z), .B(bitalign_curr_state_Z[1]), .Y(
        tap_cnt_0_sqmuxa_1_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[85]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[85]), .C(
        un10_early_flags[85]), .Y(late_flags_7_fast_Z[85]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_4 (.A(
        early_flags_pmux_126_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[43]), .D(early_flags_Z[107]), .FCI(
        early_flags_pmux_126_1_0_co0_1), .S(
        early_flags_pmux_126_1_0_wmux_4_S), .Y(
        early_flags_pmux_126_1_0_0_y5), .FCO(
        early_flags_pmux_126_1_0_co1_1));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_62 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_1_Z[32]), .Y(
        un10_early_flags[62]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[56]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[56]), .C(
        un10_early_flags[56]), .Y(late_flags_7_fast_Z[56]));
    CFG3 #( .INIT(8'h40) )  rx_err_2_sqmuxa_0_373_a2 (.A(
        restart_trng_fg_i), .B(early_flags_dec[127]), .C(
        bitalign_curr_state162_Z), .Y(N_1392));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[9]), .D(
        late_flags_Z[73]), .FCI(late_flags_pmux_126_1_1_co1_0), .S(
        late_flags_pmux_126_1_1_wmux_3_S), .Y(
        late_flags_pmux_126_1_1_y0_1), .FCO(
        late_flags_pmux_126_1_1_co0_1));
    CFG4 #( .INIT(16'h0F0E) )  emflag_cnt_1_sqmuxa_1 (.A(
        bitalign_curr_state160_Z), .B(bitalign_curr_state159_Z), .C(
        early_flags_dec[127]), .D(bitalign_curr_state161_Z), .Y(
        emflag_cnt_1_sqmuxa_1_Z));
    CFG4 #( .INIT(16'h8000) )  calc_done25_239 (.A(calc_done25_191_Z), 
        .B(calc_done25_190_Z), .C(calc_done25_189_Z), .D(
        calc_done25_188_Z), .Y(calc_done25_239_Z));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[2]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[2]), .D(GND), .FCI(
        emflag_cnt_cry_Z[1]), .S(emflag_cnt_s[2]), .Y(
        emflag_cnt_cry_Y_0[2]), .FCO(emflag_cnt_cry_Z[2]));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI6O2D1[1]  (.A(early_val_Z[1])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[1]), .Y(
        early_val_RNI6O2D1_Z[1]));
    SLE rx_BIT_ALGN_DIR (.D(un1_restart_trng_fg_6_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_BIT_ALGN_DIR_0_sqmuxa_2_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[34]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[34]), .C(
        un10_early_flags[34]), .Y(early_flags_7_fast_Z[34]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[42]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[42]), .C(
        un10_early_flags[42]), .Y(early_flags_7_fast_Z[42]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI8J6J1[2]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[2]), .D(GND), .FCI(
        timeout_cnt_cry[1]), .S(timeout_cnt_s[2]), .Y(
        timeout_cnt_RNI8J6J1_Y[2]), .FCO(timeout_cnt_cry[2]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_5_0 (
        .A(emflag_cnt_Z[5]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[5]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_4), .S(
        noearly_nolate_diff_start_7[5]), .Y(
        noearly_nolate_diff_start_7_cry_5_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[79]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[79]), .C(
        un10_early_flags[79]), .Y(late_flags_7_fast_Z[79]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[23]), 
        .D(early_flags_Z[87]), .FCI(early_flags_pmux_126_1_0_co1_5), 
        .S(early_flags_pmux_126_1_0_wmux_13_S), .Y(
        early_flags_pmux_126_1_0_y0_5), .FCO(
        early_flags_pmux_126_1_0_co0_6));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNIIHTC3[6]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[6]), .D(GND), .FCI(
        timeout_cnt_cry[5]), .S(timeout_cnt_s[6]), .Y(
        timeout_cnt_RNIIHTC3_Y[6]), .FCO(timeout_cnt_cry[6]));
    CFG2 #( .INIT(4'h1) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_0 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .Y(
        tap_cnt_0_sqmuxa_2_0));
    CFG2 #( .INIT(4'hE) )  tapcnt_final_13_m0s2 (.A(
        un1_restart_trng_fg_10_sn), .B(un1_bitalign_curr_state_12_Z), 
        .Y(tapcnt_final_13_m0s2_Z));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_0 (.A(
        early_flags_pmux_126_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[33]), .D(early_flags_Z[97]), .FCI(
        early_flags_pmux_126_1_1_co0), .S(
        early_flags_pmux_126_1_1_wmux_0_S), .Y(
        early_flags_pmux_126_1_1_y1), .FCO(
        early_flags_pmux_126_1_1_co1));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_6_0 (.A(
        emflag_cnt_Z[6]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[6]), .D(GND), .FCI(early_late_diff_8_cry_5), .S(
        early_late_diff_8[6]), .Y(early_late_diff_8_cry_6_0_Y), .FCO(
        early_late_diff_8_cry_6));
    SLE \early_flags[73]  (.D(early_flags_7_fast_Z[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[73]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_1 (.A(
        un10_tapcnt_final_1), .B(un16_tapcnt_final_1), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_0_Z), .S(
        un10_tapcnt_final_cry_1_S), .Y(un10_tapcnt_final_cry_1_Y), 
        .FCO(un10_tapcnt_final_cry_1_Z));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_108 (.A(tap_cnt_Z[4]), 
        .B(un10_early_flags_1_Z[12]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[108]));
    CFG2 #( .INIT(4'hD) )  early_late_diff_0_sqmuxa_RNIDTT8 (.A(
        early_late_diff_0_sqmuxa_1_0_Z), .B(early_late_diff_0_sqmuxa_Z)
        , .Y(early_late_diff_0_sqmuxa_1_i));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_16 (.A(
        late_flags_pmux_126_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[45]), .D(late_flags_Z[109]), .FCI(
        late_flags_pmux_126_1_1_co0_7), .S(
        late_flags_pmux_126_1_1_wmux_16_S), .Y(
        late_flags_pmux_126_1_1_y5_0), .FCO(
        late_flags_pmux_126_1_1_co1_7));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_0 (.A(
        late_flags_pmux_126_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[33]), .D(late_flags_Z[97]), .FCI(
        late_flags_pmux_126_1_1_co0), .S(
        late_flags_pmux_126_1_1_wmux_0_S), .Y(
        late_flags_pmux_126_1_1_y1), .FCO(late_flags_pmux_126_1_1_co1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[44]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[44]), .C(
        un10_early_flags[44]), .Y(late_flags_7_fast_Z[44]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_170 (.A(early_flags_Z[95]), 
        .B(early_flags_Z[94]), .C(early_flags_Z[93]), .D(
        early_flags_Z[92]), .Y(calc_done25_170_Z));
    SLE \tap_cnt[5]  (.D(N_1497_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tap_cnt_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[127]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[127]), .C(
        un10_early_flags[127]), .Y(late_flags_7_fast_Z[127]));
    CFG4 #( .INIT(16'h0BFB) )  \bitalign_curr_state_34_4_0_.m46  (.A(
        un1_retrain_adj_tap_i), .B(bitalign_curr_state13), .C(
        bitalign_curr_state_Z[0]), .D(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(N_47));
    CFG4 #( .INIT(16'hF800) )  un1_noearly_nolate_diff_start_valid (.A(
        un10_tapcnt_final_3), .B(
        un2_noearly_nolate_diff_start_validlt3), .C(
        un2_noearly_nolate_diff_start_validlto7_2_Z), .D(
        un1_early_late_diff_cry_7_Z), .Y(
        un1_noearly_nolate_diff_start_valid_Z));
    CFG4 #( .INIT(16'h0010) )  rx_trng_done1_RNO (.A(restart_trng_fg_i)
        , .B(N_1416), .C(bitalign_curr_state_Z[3]), .D(
        bitalign_curr_state_Z[2]), .Y(N_1415_i));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[71]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[71]), .C(
        un10_early_flags[71]), .Y(early_flags_7_fast_Z[71]));
    ARI1 #( .INIT(20'h5D872) )  
        \un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11[0]  (.A(tap_cnt_Z[0]), 
        .B(N_60), .C(N_89), .D(tapcnt_final_Z[0]), .FCI(GND), .S(
        un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_S[0]), .Y(
        un1_tap_cnt_0_sqmuxa_14_i_a2_RNIG1U11_Y[0]), .FCO(
        tap_cnt_17_i_m2_cry_0));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_2_sqmuxa_1_0_a2 (.A(
        tapcnt_final_upd_1_sqmuxa), .B(restart_trng_fg_i), .Y(
        tapcnt_final_upd_2_sqmuxa_1));
    CFG3 #( .INIT(8'h51) )  \bitalign_curr_state_34_4_0_.m59  (.A(
        early_flags_dec[127]), .B(late_flags_pmux), .C(
        early_flags_pmux), .Y(N_60_0));
    SLE \early_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_6 (.A(
        early_flags_pmux_126_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[57]), .D(early_flags_Z[121]), .FCI(
        early_flags_pmux_126_1_1_co0_2), .S(
        early_flags_pmux_126_1_1_wmux_6_S), .Y(
        early_flags_pmux_126_1_1_y7), .FCO(
        early_flags_pmux_126_1_1_co1_2));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_18 (.A(
        late_flags_pmux_126_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[63]), .D(late_flags_Z[127]), .FCI(
        late_flags_pmux_126_1_0_co0_8), .S(
        late_flags_pmux_126_1_0_wmux_18_S), .Y(
        late_flags_pmux_126_1_0_y7_0), .FCO(
        late_flags_pmux_126_1_0_co1_8));
    SLE \early_flags[80]  (.D(early_flags_7_fast_Z[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[80]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[25]), 
        .D(late_flags_Z[89]), .FCI(late_flags_pmux_126_1_1_co1_1), .S(
        late_flags_pmux_126_1_1_wmux_5_S), .Y(
        late_flags_pmux_126_1_1_y0_2), .FCO(
        late_flags_pmux_126_1_1_co0_2));
    SLE \late_flags[97]  (.D(late_flags_7_fast_Z[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[97]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_3_0 (
        .A(emflag_cnt_Z[3]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[3]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_2), .S(
        noearly_nolate_diff_start_7[3]), .Y(
        noearly_nolate_diff_start_7_cry_3_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_3));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI99K12[3]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[3]), .D(GND), .FCI(
        timeout_cnt_cry[2]), .S(timeout_cnt_s[3]), .Y(
        timeout_cnt_RNI99K12_Y[3]), .FCO(timeout_cnt_cry[3]));
    CFG4 #( .INIT(16'hAAAB) )  calc_done_0_sqmuxa_2_i (.A(
        restart_trng_fg_i), .B(un1_bitalign_curr_state148_8_2_Z), .C(
        early_flags_0_sqmuxa_1_Z), .D(early_flags_1_sqmuxa_1_Z), .Y(
        calc_done_0_sqmuxa_2_i_Z));
    SLE \noearly_nolate_diff_start[4]  (.D(
        noearly_nolate_diff_start_7[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_4));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_127_1_0_wmux (.A(
        emflag_cnt_Z[1]), .B(emflag_cnt_Z[0]), .C(
        late_flags_pmux_63_1_1_wmux_10_Y), .D(
        late_flags_pmux_63_1_0_wmux_10_Y), .FCI(VCC), .S(
        late_flags_pmux_127_1_0_wmux_S), .Y(late_flags_pmux_127_1_0_y0)
        , .FCO(late_flags_pmux_127_1_0_co0));
    CFG4 #( .INIT(16'h5150) )  sig_rx_BIT_ALGN_CLR_FLGS_11_iv (.A(
        restart_trng_fg_i), .B(rx_err_Z), .C(
        un1_bitalign_curr_state_1_sqmuxa_6_i_0), .D(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .Y(
        sig_rx_BIT_ALGN_CLR_FLGS_11));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_18 (.A(
        early_flags_pmux_126_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[63]), .D(early_flags_Z[127]), .FCI(
        early_flags_pmux_126_1_0_co0_8), .S(
        early_flags_pmux_126_1_0_wmux_18_S), .Y(
        early_flags_pmux_126_1_0_y7_0), .FCO(
        early_flags_pmux_126_1_0_co1_8));
    SLE \early_flags[112]  (.D(early_flags_7_fast_Z[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[112]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_12 (.A(
        late_flags_pmux_126_1_1_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[37]), .D(late_flags_Z[101]), .FCI(
        late_flags_pmux_126_1_1_co0_5), .S(
        late_flags_pmux_126_1_1_wmux_12_S), .Y(
        late_flags_pmux_126_1_1_y1_0), .FCO(
        late_flags_pmux_126_1_1_co1_5));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[4]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[4]), .D(GND), .FCI(
        emflag_cnt_cry_Z[3]), .S(emflag_cnt_s[4]), .Y(
        emflag_cnt_cry_Y_0[4]), .FCO(emflag_cnt_cry_Z[4]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[8]), 
        .D(early_flags_Z[72]), .FCI(early_flags_pmux_63_1_1_co1_0), .S(
        early_flags_pmux_63_1_1_wmux_3_S), .Y(
        early_flags_pmux_63_1_1_y0_1), .FCO(
        early_flags_pmux_63_1_1_co0_1));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_14 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[3]), .C(un10_early_flags_1_Z[6]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[14]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_41 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_0[40]), .C(
        un10_early_flags_2_Z[37]), .Y(un10_early_flags[41]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[5]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[5]), .D(GND), .FCI(
        emflag_cnt_cry_Z[4]), .S(emflag_cnt_s[5]), .Y(
        emflag_cnt_cry_Y_0[5]), .FCO(emflag_cnt_cry_Z[5]));
    CFG4 #( .INIT(16'h0D00) )  calc_done27 (.A(un34), .B(
        un16_tapcnt_final_cry_7_Z), .C(calc_done25_Z), .D(
        un1_noearly_nolate_diff_start_valid_Z), .Y(calc_done27_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[76]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[76]), .C(
        un10_early_flags[76]), .Y(late_flags_7_fast_Z[76]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_16 (.A(
        late_flags_pmux_63_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[44]), .D(late_flags_Z[108]), .FCI(
        late_flags_pmux_63_1_1_co0_7), .S(
        late_flags_pmux_63_1_1_wmux_16_S), .Y(
        late_flags_pmux_63_1_1_y5_0), .FCO(
        late_flags_pmux_63_1_1_co1_7));
    SLE \late_flags[58]  (.D(late_flags_7_fast_Z[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[58]));
    SLE \late_flags[108]  (.D(late_flags_7_fast_Z[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[108]));
    CFG3 #( .INIT(8'hDC) )  un1_early_flags_1_sqmuxa_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(early_flags_1_sqmuxa_Z), .C(
        bitalign_curr_state156_Z), .Y(un1_early_flags_1_sqmuxa_1_Z));
    SLE \early_flags[18]  (.D(early_flags_7_fast_Z[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[18]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[111]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[111]), .C(
        un10_early_flags[111]), .Y(late_flags_7_fast_Z[111]));
    SLE \rst_cnt[1]  (.D(rst_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[1]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_110 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[64]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_1_Z[40]), .Y(
        un10_early_flags[110]));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state148_5_4 (.A(
        bitalign_curr_state154_3_Z), .B(bitalign_curr_state149_Z), .C(
        bitalign_curr_state148_Z), .Y(un1_bitalign_curr_state148_5_4_Z)
        );
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_10 (.A(
        early_flags_pmux_63_1_1_y21), .B(early_flags_pmux_63_1_1_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_63_1_1_co0_4), .S(
        early_flags_pmux_63_1_1_wmux_10_S), .Y(
        early_flags_pmux_63_1_1_wmux_10_Y), .FCO(
        early_flags_pmux_63_1_1_co1_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[100]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[100]), .C(
        un10_early_flags[100]), .Y(early_flags_7_fast_Z[100]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_55 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_47_0_Z), .Y(
        un10_early_flags[55]));
    SLE \early_flags[90]  (.D(early_flags_7_fast_Z[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[90]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_128 (.A(late_flags_Z[119]), 
        .B(late_flags_Z[118]), .C(late_flags_Z[117]), .D(
        late_flags_Z[116]), .Y(calc_done25_128_Z));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_1_wmux_8 (.A(
        late_flags_pmux_63_1_1_y0_3), .B(late_flags_pmux_63_1_1_y3), 
        .C(late_flags_pmux_63_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co0_3), .S(
        late_flags_pmux_63_1_1_wmux_8_S), .Y(late_flags_pmux_63_1_1_y9)
        , .FCO(late_flags_pmux_63_1_1_co1_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[10]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[10]), .C(
        un10_early_flags[10]), .Y(late_flags_7_fast_Z[10]));
    ARI1 #( .INIT(20'h40D00) )  \emflag_cnt_cry_cy[0]  (.A(VCC), .B(
        N_1456_1), .C(bitalign_curr_state_Z[1]), .D(
        un1_restart_trng_fg_9_0_443_0), .FCI(VCC), .S(
        emflag_cnt_cry_cy_S_0[0]), .Y(emflag_cnt_cry_cy_Y_0[0]), .FCO(
        emflag_cnt_cry_cy));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[87]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[87]), .C(
        un10_early_flags[87]), .Y(late_flags_7_fast_Z[87]));
    SLE \late_flags[83]  (.D(late_flags_7_fast_Z[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[83]));
    SLE \early_flags[82]  (.D(early_flags_7_fast_Z[82]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[82]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_87 (.A(
        un10_early_flags_1_Z[20]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_3_Z[87]), .Y(
        un10_early_flags[87]));
    SLE \wait_cnt[0]  (.D(wait_cnt_4_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(wait_cnt_Z[0]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_0 (.A(
        un16_tapcnt_final_0), .B(un10_tapcnt_final_0), .C(GND), .D(GND)
        , .FCI(GND), .S(un16_tapcnt_final_cry_0_S), .Y(
        un16_tapcnt_final_cry_0_Y), .FCO(un16_tapcnt_final_cry_0_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[57]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[57]), .C(
        un10_early_flags[57]), .Y(early_flags_7_fast_Z[57]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_4 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_2_0[0]), .D(
        un10_early_flags_2_Z[4]), .Y(un10_early_flags[4]));
    SLE \no_early_no_late_val_st1[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[6]));
    SLE \late_flags[68]  (.D(late_flags_7_fast_Z[68]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[68]));
    CFG2 #( .INIT(4'h1) )  \bitalign_curr_state_34_4_0_.m8  (.A(
        bitalign_curr_state_Z[0]), .B(BIT_ALGN_OOR_c), .Y(N_9));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_65 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[6]), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[65]));
    CFG3 #( .INIT(8'h80) )  early_late_diff_0_sqmuxa (.A(
        late_flags_pmux), .B(late_last_set15_Z), .C(
        bitalign_curr_state161_Z), .Y(early_late_diff_0_sqmuxa_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_40 (.A(
        un10_early_flags_2_0[40]), .B(un10_early_flags_1_Z[0]), .C(
        un10_early_flags_1_Z[40]), .Y(un10_early_flags[40]));
    CFG4 #( .INIT(16'hFFFE) )  early_last_set_0_sqmuxa_i (.A(
        un1_restart_trng_fg_10_sn_1), .B(early_last_set_1_sqmuxa_1_3_Z)
        , .C(early_val_0_sqmuxa_1_0_Z), .D(tap_cnt_0_sqmuxa_1_Z), .Y(
        early_last_set_0_sqmuxa_i_Z));
    SLE \early_late_diff[4]  (.D(early_late_diff_8[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[4]));
    CFG4 #( .INIT(16'hFF3B) )  un1_bitalign_curr_state_16_1 (.A(
        bitalign_curr_state_Z[2]), .B(N_117_mux_1), .C(
        bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[4]), .Y(
        un1_bitalign_curr_state_16_1_Z));
    SLE \late_flags[13]  (.D(late_flags_7_fast_Z[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[13]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_0_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_126_1_0_co1_3), .S(
        late_flags_pmux_126_1_0_wmux_9_S), .Y(
        late_flags_pmux_126_1_0_wmux_9_Y), .FCO(
        late_flags_pmux_126_1_0_co0_4));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[95]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[95]), .C(
        un10_early_flags[95]), .Y(late_flags_7_fast_Z[95]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_47_0 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[6]), .Y(un10_early_flags_47_0_Z));
    SLE \timeout_cnt[6]  (.D(timeout_cnt_s[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[6]));
    SLE \tap_cnt[1]  (.D(N_30_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[1]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_2 (.A(
        late_flags_pmux_63_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[50]), .D(late_flags_Z[114]), .FCI(
        late_flags_pmux_63_1_0_co0_0), .S(
        late_flags_pmux_63_1_0_wmux_2_S), .Y(
        late_flags_pmux_63_1_0_0_y3), .FCO(
        late_flags_pmux_63_1_0_co1_0));
    CFG3 #( .INIT(8'h20) )  \bitalign_curr_state_34_4_0_.m66_2  (.A(
        bitalign_curr_state_Z[3]), .B(bitalign_curr_state_Z[4]), .C(
        N_65), .Y(m66_1));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[6]  (.A(
        no_early_no_late_val_end1_Z[6]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[6]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[20]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[20]), .C(
        un10_early_flags[20]), .Y(early_flags_7_fast_Z[20]));
    SLE \early_flags[3]  (.D(early_flags_7_fast_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[3]));
    CFG4 #( .INIT(16'hFF9C) )  \wait_cnt_4[1]  (.A(wait_cnt_Z[0]), .B(
        wait_cnt_Z[1]), .C(bitalign_curr_state152_3_Z), .D(
        un1_restart_trng_fg_Z), .Y(wait_cnt_4_Z[1]));
    CFG2 #( .INIT(4'hD) )  early_val_0_sqmuxa_1_i (.A(
        early_cur_set_0_sqmuxa_1_Z), .B(un1_tap_cnt_0_sqmuxa_6_0), .Y(
        early_val_0_sqmuxa_1_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[80]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[80]), .C(
        un10_early_flags[80]), .Y(early_flags_7_fast_Z[80]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_100 (.A(
        un10_early_flags_1_Z[36]), .B(un10_early_flags_1_Z[64]), .C(
        un10_early_flags_2_0[100]), .Y(un10_early_flags[100]));
    CFG2 #( .INIT(4'h8) )  sig_rx_BIT_ALGN_CLR_FLGS14 (.A(CO0_0), .B(
        cnt_Z[1]), .Y(sig_rx_BIT_ALGN_CLR_FLGS14_Z));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_0_0 (.A(
        emflag_cnt_Z[0]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[0]), .D(GND), .FCI(early_late_diff_8_cry_0_0_cy_Z), 
        .S(early_late_diff_8[0]), .Y(early_late_diff_8_cry_0_0_Y), 
        .FCO(early_late_diff_8_cry_0));
    CFG4 #( .INIT(16'h8000) )  early_flags_dec_127 (.A(emflag_cnt_Z[2])
        , .B(early_flags_dec_127_4_Z), .C(emflag_cnt_Z[1]), .D(
        emflag_cnt_Z[0]), .Y(early_flags_dec[127]));
    SLE \late_flags[54]  (.D(late_flags_7_fast_Z[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[54]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_2 (.A(
        early_flags_pmux_126_1_1_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[49]), .D(early_flags_Z[113]), .FCI(
        early_flags_pmux_126_1_1_co0_0), .S(
        early_flags_pmux_126_1_1_wmux_2_S), .Y(
        early_flags_pmux_126_1_1_y3), .FCO(
        early_flags_pmux_126_1_1_co1_0));
    SLE \late_flags[43]  (.D(late_flags_7_fast_Z[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[43]));
    SLE \early_flags[92]  (.D(early_flags_7_fast_Z[92]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[92]));
    CFG3 #( .INIT(8'h08) )  bitalign_curr_state_1_sqmuxa_4 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state149_Z), 
        .C(BIT_ALGN_ERR_0_c), .Y(bitalign_curr_state_1_sqmuxa_4_Z));
    SLE \early_flags[124]  (.D(early_flags_7_fast_Z[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[124]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[47]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[47]), .C(
        un10_early_flags[47]), .Y(early_flags_7_fast_Z[47]));
    CFG2 #( .INIT(4'h4) )  bitalign_curr_state89 (.A(early_flags_pmux), 
        .B(late_flags_pmux), .Y(bitalign_curr_state89_Z));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_0_wmux_20 (.A(
        late_flags_pmux_63_1_0_y0_8), .B(late_flags_pmux_63_1_0_y3_0), 
        .C(late_flags_pmux_63_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co0_9), .S(
        late_flags_pmux_63_1_0_wmux_20_S), .Y(
        late_flags_pmux_63_1_0_0_y21), .FCO(
        late_flags_pmux_63_1_0_co1_9));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[15]), 
        .D(late_flags_Z[79]), .FCI(late_flags_pmux_126_1_0_co1_6), .S(
        late_flags_pmux_126_1_0_wmux_15_S), .Y(
        late_flags_pmux_126_1_0_y0_6), .FCO(
        late_flags_pmux_126_1_0_co0_7));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[60]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[60]), .C(
        un10_early_flags[60]), .Y(early_flags_7_fast_Z[60]));
    CFG2 #( .INIT(4'h6) )  \cnt_RNO[1]  (.A(CO0_0), .B(cnt_Z[1]), .Y(
        cnt_RNO_Z[1]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_225 (.A(calc_done25_135_Z), 
        .B(calc_done25_134_Z), .C(calc_done25_133_Z), .D(
        calc_done25_132_Z), .Y(calc_done25_225_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_86 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[6]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[6]), .Y(
        un10_early_flags[86]));
    SLE \early_flags[45]  (.D(early_flags_7_fast_Z[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[45]));
    CFG3 #( .INIT(8'h46) )  \bitalign_curr_state_34_4_0_.m12  (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state_Z[0]), 
        .C(bitalign_curr_state61), .Y(N_114_mux));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_100_2_0 (.A(
        un10_early_flags_2_Z[4]), .B(tap_cnt_Z[4]), .Y(
        un10_early_flags_2_0[100]));
    SLE \late_flags[122]  (.D(late_flags_7_fast_Z[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[122]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_16_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[3]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[16]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_58 (.A(tap_cnt_Z[6]), 
        .B(un10_early_flags_1_Z[10]), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[58]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[62]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[62]), .C(
        un10_early_flags[62]), .Y(late_flags_7_fast_Z[62]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_157 (.A(late_flags_Z[3]), 
        .B(late_flags_Z[2]), .C(late_flags_Z[1]), .D(late_flags_Z[0]), 
        .Y(calc_done25_157_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_18 (.A(
        late_flags_pmux_63_1_0_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[62]), .D(late_flags_Z[126]), .FCI(
        late_flags_pmux_63_1_0_co0_8), .S(
        late_flags_pmux_63_1_0_wmux_18_S), .Y(
        late_flags_pmux_63_1_0_y7_0), .FCO(
        late_flags_pmux_63_1_0_co1_8));
    CFG3 #( .INIT(8'hB1) )  \bitalign_curr_state_34_4_0_.m13  (.A(
        bitalign_curr_state_Z[1]), .B(N_11), .C(N_114_mux), .Y(N_14));
    CFG4 #( .INIT(16'h0040) )  bitalign_curr_state164 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state152_1_Z), .D(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state164_Z));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[1]  (.A(N_79), .B(N_63_0), .Y(
        N_30_i));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_24_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[2]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[24]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_19 (.A(
        early_flags_pmux_63_1_1_y7_0), .B(early_flags_pmux_63_1_1_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co1_8), .S(
        early_flags_pmux_63_1_1_wmux_19_S), .Y(
        early_flags_pmux_63_1_1_y0_8), .FCO(
        early_flags_pmux_63_1_1_co0_9));
    SLE \late_flags[22]  (.D(late_flags_7_fast_Z[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[22]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_161 (.A(early_flags_Z[115]), 
        .B(early_flags_Z[114]), .C(early_flags_Z[113]), .D(
        early_flags_Z[112]), .Y(calc_done25_161_Z));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_7 (.A(
        un16_tapcnt_final_7), .B(un10_tapcnt_final_7), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_6_Z), .S(
        un16_tapcnt_final_cry_7_S), .Y(un16_tapcnt_final_cry_7_Y), 
        .FCO(un16_tapcnt_final_cry_7_Z));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[2]  (.A(
        no_early_no_late_val_end1_Z[2]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[2]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[2]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_3 (.A(
        un10_tapcnt_final_3), .B(un16_tapcnt_final_3), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_2_Z), .S(
        un10_tapcnt_final_cry_3_S), .Y(un10_tapcnt_final_cry_3_Y), 
        .FCO(un10_tapcnt_final_cry_3_Z));
    CFG4 #( .INIT(16'h0400) )  un10_early_flags_79 (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[6]), .C(tap_cnt_Z[5]), .D(
        un10_early_flags_1_0[15]), .Y(un10_early_flags[79]));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.m43_0_a2_0  (
        .A(BIT_ALGN_ERR_0_c), .B(retrain_reg_Z[2]), .Y(
        un1_rx_BIT_ALGN_START));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[1]  (.A(
        no_early_no_late_val_end1_Z[1]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[1]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[1]));
    CFG2 #( .INIT(4'hE) )  rx_err_1_sqmuxa_RNIG5FO1 (.A(
        rx_err_1_sqmuxa_Z), .B(emflag_cntlde_4), .Y(emflag_cnte));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_4 (.A(
        late_flags_pmux_126_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[43]), .D(late_flags_Z[107]), .FCI(
        late_flags_pmux_126_1_0_co0_1), .S(
        late_flags_pmux_126_1_0_wmux_4_S), .Y(
        late_flags_pmux_126_1_0_0_y5), .FCO(
        late_flags_pmux_126_1_0_co1_1));
    CFG4 #( .INIT(16'h72AA) )  \bitalign_curr_state_34_4_0_.m30  (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state41_Z), .C(
        bit_align_dly_done_Z), .D(bitalign_curr_state_Z[1]), .Y(N_31));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[23]), 
        .D(late_flags_Z[87]), .FCI(late_flags_pmux_126_1_0_co1_5), .S(
        late_flags_pmux_126_1_0_wmux_13_S), .Y(
        late_flags_pmux_126_1_0_y0_5), .FCO(
        late_flags_pmux_126_1_0_co0_6));
    CFG4 #( .INIT(16'h0001) )  calc_done25_190 (.A(early_flags_Z[15]), 
        .B(early_flags_Z[14]), .C(early_flags_Z[13]), .D(
        early_flags_Z[12]), .Y(calc_done25_190_Z));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_68 (.A(tap_cnt_Z[2]), 
        .B(tap_cnt_Z[6]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[68]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_14 (.A(
        late_flags_pmux_63_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[52]), .D(late_flags_Z[116]), .FCI(
        late_flags_pmux_63_1_1_co0_6), .S(
        late_flags_pmux_63_1_1_wmux_14_S), .Y(
        late_flags_pmux_63_1_1_y3_0), .FCO(
        late_flags_pmux_63_1_1_co1_6));
    SLE \late_flags[64]  (.D(late_flags_7_fast_Z[64]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[64]));
    CFG2 #( .INIT(4'h8) )  bitalign_curr_state155_1 (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state155_1_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[7]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[7]), .C(
        un10_early_flags[7]), .Y(early_flags_7_fast_Z[7]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[24]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[24]), .C(
        un10_early_flags[24]), .Y(early_flags_7_fast_Z[24]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[84]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[84]), .C(
        un10_early_flags[84]), .Y(early_flags_7_fast_Z[84]));
    SLE \no_early_no_late_val_st1[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[59]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[59]), .C(
        un10_early_flags[59]), .Y(early_flags_7_fast_Z[59]));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_3_sqmuxa_1_0_a2 (.A(
        tapcnt_final_upd_2_sqmuxa), .B(restart_trng_fg_i), .Y(
        tapcnt_final_upd_3_sqmuxa_1));
    CFG4 #( .INIT(16'hFFF8) )  un1_bitalign_curr_state_1_sqmuxa_2 (.A(
        tap_cnt_0_sqmuxa_1_0_Z), .B(tap_cnt_0_sqmuxa_2_0), .C(
        bitalign_curr_state_1_sqmuxa_4_Z), .D(tap_cnt_0_sqmuxa_1_Z), 
        .Y(un1_bitalign_curr_state_1_sqmuxa_2_i_0));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNIF13D1[4]  (.A(early_val_Z[4])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[4]), .Y(
        early_val_RNIF13D1_Z[4]));
    CFG3 #( .INIT(8'h40) )  un10_early_flags_17 (.A(N_1498), .B(
        un10_early_flags_2_Z[8]), .C(un10_early_flags_2_0[16]), .Y(
        un10_early_flags[17]));
    SLE \late_flags[72]  (.D(late_flags_7_fast_Z[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[72]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_0 (.A(
        early_flags_pmux_63_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[32]), .D(early_flags_Z[96]), .FCI(
        early_flags_pmux_63_1_1_co0), .S(
        early_flags_pmux_63_1_1_wmux_0_S), .Y(
        early_flags_pmux_63_1_1_y1), .FCO(early_flags_pmux_63_1_1_co1));
    SLE \timeout_cnt[0]  (.D(timeout_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[0]));
    SLE \late_flags[114]  (.D(late_flags_7_fast_Z[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[114]));
    SLE \late_flags[3]  (.D(late_flags_7_fast_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[3]));
    SLE \late_flags[100]  (.D(late_flags_7_fast_Z[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[100]));
    CFG4 #( .INIT(16'h4000) )  bit_align_dly_done_0_sqmuxa (.A(
        bitalign_curr_state_Z[4]), .B(rx_trng_done_Z), .C(
        bitalign_curr_state161_2_Z), .D(bitalign_curr_state159_2_Z), 
        .Y(bit_align_dly_done_0_sqmuxa_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[18]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[18]), .C(
        un10_early_flags[18]), .Y(late_flags_7_fast_Z[18]));
    CFG4 #( .INIT(16'hDDEC) )  \bitalign_curr_state_34_4_0_.m91  (.A(
        bitalign_curr_state_Z[2]), .B(m91_1), .C(N_116_mux), .D(
        m91_1_0), .Y(N_92));
    CFG4 #( .INIT(16'hFEFC) )  mv_dn_fg_0_sqmuxa_i_o2 (.A(
        bitalign_curr_state148_Z), .B(bitalign_curr_state_1_sqmuxa_4_Z)
        , .C(restart_trng_fg_i), .D(N_61), .Y(mv_dn_fg_0_sqmuxa_i_o2_Z)
        );
    CFG4 #( .INIT(16'hFDFC) )  un1_restart_trng_fg_8 (.A(
        early_flags_pmux), .B(un1_tap_cnt_0_sqmuxa_6_0), .C(
        restart_trng_fg_i), .D(early_val_0_sqmuxa_1_0_Z), .Y(
        un1_restart_trng_fg_8_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[64]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[64]), .C(
        un10_early_flags[64]), .Y(early_flags_7_fast_Z[64]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_155 (.A(late_flags_Z[27]), 
        .B(late_flags_Z[26]), .C(late_flags_Z[25]), .D(
        late_flags_Z[24]), .Y(calc_done25_155_Z));
    SLE \late_flags[93]  (.D(late_flags_7_fast_Z[93]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[93]));
    SLE \late_flags[89]  (.D(late_flags_7_fast_Z[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[89]));
    CFG4 #( .INIT(16'hFFFE) )  late_cur_set_0_sqmuxa_i (.A(
        un1_restart_trng_fg_10_sn_1), .B(tap_cnt_0_sqmuxa_1_Z), .C(
        early_last_set_1_sqmuxa_1_3_Z), .D(
        un1_bitalign_curr_state_2_sqmuxa_Z), .Y(
        late_cur_set_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[38]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[38]), .C(
        un10_early_flags[38]), .Y(early_flags_7_fast_Z[38]));
    ARI1 #( .INIT(20'h574B8) )  \tapcnt_final_RNISU155[4]  (.A(
        tap_cnt_Z[4]), .B(un1_tap_cnt_0_sqmuxa_14_0_Z[1]), .C(N_60), 
        .D(tapcnt_final_Z[4]), .FCI(tap_cnt_17_i_m2_cry_3), .S(N_76), 
        .Y(tapcnt_final_RNISU155_Y[4]), .FCO(tap_cnt_17_i_m2_cry_4));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[123]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[123]), .C(
        un10_early_flags[123]), .Y(early_flags_7_fast_Z[123]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_32_2_0 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[32]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[97]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[97]), .C(
        un10_early_flags[97]), .Y(late_flags_7_fast_Z[97]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_51 (.A(
        un10_early_flags_1_Z[3]), .B(un10_early_flags_2_0[48]), .C(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[51]));
    SLE \late_flags[32]  (.D(late_flags_7_fast_Z[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[32]));
    CFG2 #( .INIT(4'hE) )  un1_bitalign_curr_state_15_1 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[4]), .Y(
        un1_bitalign_curr_state_15_1_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[8]  (.A(VCC), .B(
        rst_cnt_Z[8]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[7]), .S(
        rst_cnt_s[8]), .Y(rst_cnt_cry_Y_0[8]), .FCO(rst_cnt_cry_Z[8]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_7 (.A(
        late_flags_pmux_63_1_0_0_y7), .B(late_flags_pmux_63_1_0_0_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co1_2), .S(
        late_flags_pmux_63_1_0_wmux_7_S), .Y(
        late_flags_pmux_63_1_0_y0_3), .FCO(
        late_flags_pmux_63_1_0_co0_3));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[16]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[16]), .C(
        un10_early_flags[16]), .Y(early_flags_7_fast_Z[16]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[35]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[35]), .C(
        un10_early_flags[35]), .Y(early_flags_7_fast_Z[35]));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_10_2 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[10]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_0 (.A(late_val_Z[0])
        , .B(early_val_Z[0]), .C(GND), .D(GND), .FCI(GND), .S(
        tapcnt_final27_cry_0_S), .Y(tapcnt_final27_cry_0_Y), .FCO(
        tapcnt_final27_cry_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[80]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[80]), .C(
        un10_early_flags[80]), .Y(late_flags_7_fast_Z[80]));
    SLE \late_flags[119]  (.D(late_flags_7_fast_Z[119]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[119]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_67_2 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[67]));
    CFG4 #( .INIT(16'h8000) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(tap_cnt_0_sqmuxa_2_0), .C(
        bitalign_curr_state_Z[1]), .D(un1_bitalign_curr_state151_Z), 
        .Y(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_Z));
    SLE \late_flags[9]  (.D(late_flags_7_fast_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[9]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[5]  (.A(
        tapcnt_final_Z[5]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[5]), .Y(
        tapcnt_final_13_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[6]), 
        .D(early_flags_Z[70]), .FCI(early_flags_pmux_63_1_0_co1_4), .S(
        early_flags_pmux_63_1_0_wmux_11_S), .Y(
        early_flags_pmux_63_1_0_y0_4), .FCO(
        early_flags_pmux_63_1_0_co0_5));
    SLE \late_flags[19]  (.D(late_flags_7_fast_Z[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[19]));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_6 (.A(
        tapcnt_final_upd_Z[6]), .B(tapcnt_final_Z[6]), .C(tap_cnt_Z[6])
        , .D(N_1416), .Y(bitalign_curr_state61_6_Z));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[3]  (.A(
        no_early_no_late_val_end1_Z[3]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[3]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[3]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNI1B921[4]  (.A(
        no_early_no_late_val_st1_Z[4]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[4]), .Y(
        un1_no_early_no_late_val_st1_1_1[4]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_72_2_0 (.A(tap_cnt_Z[2]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[5]), .Y(
        un10_early_flags_2_0[72]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_61 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_2_Z[37]), .Y(
        un10_early_flags[61]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_19 (.A(
        late_flags_pmux_126_1_1_y7_0), .B(late_flags_pmux_126_1_1_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co1_8), .S(
        late_flags_pmux_126_1_1_wmux_19_S), .Y(
        late_flags_pmux_126_1_1_y0_8), .FCO(
        late_flags_pmux_126_1_1_co0_9));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[28]), 
        .D(late_flags_Z[92]), .FCI(late_flags_pmux_63_1_1_co1_7), .S(
        late_flags_pmux_63_1_1_wmux_17_S), .Y(
        late_flags_pmux_63_1_1_y0_7), .FCO(
        late_flags_pmux_63_1_1_co0_8));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_16 (.A(
        un10_early_flags_1_Z[16]), .B(un10_early_flags_2_Z[8]), .C(
        un10_early_flags_2_0[16]), .Y(un10_early_flags[16]));
    CFG4 #( .INIT(16'h1F0E) )  \bitalign_curr_state_34_4_0_.m50  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        m50_1_1), .D(N_47), .Y(N_51));
    SLE \early_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[1]));
    CFG4 #( .INIT(16'hFFFE) )  un2_noearly_nolate_diff_nxt_validlto7_2 
        (.A(un16_tapcnt_final_7), .B(un16_tapcnt_final_6), .C(
        un16_tapcnt_final_5), .D(un16_tapcnt_final_4), .Y(
        un2_noearly_nolate_diff_nxt_validlto7_2_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[2]  (.A(VCC), .B(
        rst_cnt_Z[2]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[1]), .S(
        rst_cnt_s[2]), .Y(rst_cnt_cry_Y_0[2]), .FCO(rst_cnt_cry_Z[2]));
    SLE \early_flags[24]  (.D(early_flags_7_fast_Z[24]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[24]));
    SLE \late_flags[49]  (.D(late_flags_RNO_Z[49]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[49]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_141 (.A(late_flags_Z[67]), 
        .B(late_flags_Z[66]), .C(late_flags_Z[65]), .D(
        late_flags_Z[64]), .Y(calc_done25_141_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[13]), 
        .D(late_flags_Z[77]), .FCI(late_flags_pmux_126_1_1_co1_6), .S(
        late_flags_pmux_126_1_1_wmux_15_S), .Y(
        late_flags_pmux_126_1_1_y0_6), .FCO(
        late_flags_pmux_126_1_1_co0_7));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_124 (.A(
        un10_early_flags_1_Z[12]), .B(tap_cnt_Z[1]), .C(
        un10_early_flags_1_Z[48]), .D(un10_early_flags_1_Z[64]), .Y(
        un10_early_flags[124]));
    CFG3 #( .INIT(8'hE0) )  \wait_cnt_4_RNO[2]  (.A(wait_cnt_Z[1]), .B(
        wait_cnt_Z[0]), .C(bitalign_curr_state152_3_Z), .Y(CO1));
    CFG4 #( .INIT(16'h0001) )  bitalign_curr_state61_0_0_RNIQOA01 (.A(
        bitalign_curr_state61_0), .B(bitalign_curr_state61_NE_4_Z), .C(
        bitalign_curr_state61_5_Z), .D(bitalign_curr_state61_4_Z), .Y(
        bitalign_curr_state61));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_4_2 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[4]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_127_1_0_wmux_0 (.A(
        early_flags_pmux_127_1_0_y0), .B(emflag_cnt_Z[0]), .C(
        early_flags_pmux_126_1_1_wmux_10_Y), .D(
        early_flags_pmux_126_1_0_wmux_10_Y), .FCI(
        early_flags_pmux_127_1_0_co0), .S(
        early_flags_pmux_127_1_0_wmux_0_S), .Y(early_flags_pmux), .FCO(
        early_flags_pmux_127_1_0_co1));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_5 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_2_Z[4]), .Y(un10_early_flags[5]));
    SLE \early_flags[116]  (.D(early_flags_7_fast_Z[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[116]));
    CFG2 #( .INIT(4'h1) )  \bitalign_curr_state_34_4_0_.m98_1  (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[1]), .Y(
        N_117_mux_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[8]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[8]), .C(
        un10_early_flags[8]), .Y(early_flags_7_fast_Z[8]));
    CFG3 #( .INIT(8'h1D) )  \tapcnt_final_13_RNO_1[6]  (.A(
        no_early_no_late_val_st1_Z[6]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[6]), .Y(
        un1_no_early_no_late_val_st1_1_1[6]));
    SLE \no_early_no_late_val_st2[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[6]));
    CFG4 #( .INIT(16'hEDDE) )  \wait_cnt_4[2]  (.A(wait_cnt_Z[2]), .B(
        un1_restart_trng_fg_Z), .C(bitalign_curr_state152_3_Z), .D(CO1)
        , .Y(wait_cnt_4_Z[2]));
    ARI1 #( .INIT(20'h51045) )  tapcnt_final_upd_8_cry_4_0 (.A(
        tap_cnt_Z[4]), .B(mv_dn_fg_0_sqmuxa_i_o2_Z), .C(mv_up_fg_Z), 
        .D(N_100), .FCI(tapcnt_final_upd_8_cry_3), .S(
        tapcnt_final_upd_8[4]), .Y(tapcnt_final_upd_8_cry_4_0_Y), .FCO(
        tapcnt_final_upd_8_cry_4));
    SLE \emflag_cnt[5]  (.D(emflag_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[5]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_0_wmux_8 (.A(
        late_flags_pmux_126_1_0_y0_3), .B(late_flags_pmux_126_1_0_0_y3)
        , .C(late_flags_pmux_126_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co0_3), .S(
        late_flags_pmux_126_1_0_wmux_8_S), .Y(
        late_flags_pmux_126_1_0_0_y9), .FCO(
        late_flags_pmux_126_1_0_co1_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[64]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[64]), .C(
        un10_early_flags[64]), .Y(late_flags_7_fast_Z[64]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_181 (.A(early_flags_Z[35]), 
        .B(early_flags_Z[34]), .C(early_flags_Z[33]), .D(
        early_flags_Z[32]), .Y(calc_done25_181_Z));
    CFG3 #( .INIT(8'hC8) )  un1_bitalign_curr_state_2_sqmuxa (.A(
        emflag_cnt_0_sqmuxa), .B(bitalign_curr_state89_Z), .C(
        bitalign_curr_state159_Z), .Y(
        un1_bitalign_curr_state_2_sqmuxa_Z));
    CFG3 #( .INIT(8'hCD) )  \bitalign_curr_state_34_4_0_.m37  (.A(
        m37_1_1), .B(m37), .C(early_flags_dec[127]), .Y(i12_mux_0));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_44 (.A(
        un10_early_flags_2_0[44]), .B(un10_early_flags_1_Z[32]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[44]));
    SLE \early_flags[13]  (.D(early_flags_7_fast_Z[13]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[13]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_6 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_2_0[0]), .C(
        un10_early_flags_2_Z[6]), .Y(un10_early_flags[6]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[14]), 
        .D(late_flags_Z[78]), .FCI(late_flags_pmux_63_1_0_co1_6), .S(
        late_flags_pmux_63_1_0_wmux_15_S), .Y(
        late_flags_pmux_63_1_0_y0_6), .FCO(
        late_flags_pmux_63_1_0_co0_7));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[90]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[90]), .C(
        un10_early_flags[90]), .Y(early_flags_7_fast_Z[90]));
    CFG4 #( .INIT(16'hA0A3) )  \bitalign_curr_state_34_4_0_.m7  (.A(
        m7_1_1), .B(bitalign_curr_state12_Z), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        N_8));
    SLE \tap_cnt[4]  (.D(N_24_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[4]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_131 (.A(late_flags_Z[123]), 
        .B(late_flags_Z[122]), .C(late_flags_Z[121]), .D(
        late_flags_Z[120]), .Y(calc_done25_131_Z));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_60 (.A(tap_cnt_Z[6]), 
        .B(un10_early_flags_1_Z[12]), .C(un10_early_flags_1_Z[0]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[60]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_168 (.A(early_flags_Z[87]), 
        .B(early_flags_Z[86]), .C(early_flags_Z[85]), .D(
        early_flags_Z[84]), .Y(calc_done25_168_Z));
    SLE \early_flags[26]  (.D(early_flags_7_fast_Z[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[26]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_93 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_1_Z[24]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[69]), .Y(
        un10_early_flags[93]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_10_1 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_1_Z[10]));
    SLE \early_flags[27]  (.D(early_flags_7_fast_Z[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[27]));
    CFG4 #( .INIT(16'h0015) )  early_cur_set_0_sqmuxa_1 (.A(
        restart_trng_fg_i), .B(un1_early_last_set_1_sqmuxa_1_1_tz_Z), 
        .C(early_flags_pmux), .D(early_last_set_1_sqmuxa_1_3_Z), .Y(
        early_cur_set_0_sqmuxa_1_Z));
    SLE \late_flags[115]  (.D(late_flags_7_fast_Z[115]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[115]));
    CFG2 #( .INIT(4'h4) )  \tapcnt_final_upd_8[1]  (.A(
        mv_dn_fg_0_sqmuxa_i_o2_Z), .B(tap_cnt_Z[1]), .Y(
        tapcnt_final_upd_8_Z[1]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_52_2_0 (.A(
        un10_early_flags_2_Z[4]), .B(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[52]));
    SLE \tap_cnt[3]  (.D(N_26_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[3]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[19]), 
        .D(late_flags_Z[83]), .FCI(late_flags_pmux_126_1_0_0_co1), .S(
        late_flags_pmux_126_1_0_wmux_1_S), .Y(
        late_flags_pmux_126_1_0_y0_0), .FCO(
        late_flags_pmux_126_1_0_co0_0));
    SLE \early_flags[59]  (.D(early_flags_7_fast_Z[59]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[59]));
    CFG2 #( .INIT(4'h1) )  bitalign_curr_state161_2 (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state161_2_Z));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_69_2 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[69]));
    SLE \timeout_cnt[2]  (.D(timeout_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[2]));
    SLE \no_early_no_late_val_end1[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[5]));
    CFG2 #( .INIT(4'h2) )  early_flags_1_sqmuxa_1 (.A(
        bitalign_curr_state148_Z), .B(bitalign_curr_state12_Z), .Y(
        early_flags_1_sqmuxa_1_Z));
    SLE \early_flags[21]  (.D(early_flags_7_fast_Z[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[21]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[1]  (.A(
        tapcnt_final_Z[1]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[1]), .Y(
        tapcnt_final_13_Z[1]));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_nxt_8_cry_0_0_cy (
        .A(VCC), .B(un1_restart_trng_fg_5_Z), .C(GND), .D(GND), .FCI(
        VCC), .S(noearly_nolate_diff_nxt_8_cry_0_0_cy_S), .Y(
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_19 (.A(
        early_flags_pmux_63_1_0_y7_0), .B(early_flags_pmux_63_1_0_y5_0)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co1_8), .S(
        early_flags_pmux_63_1_0_wmux_19_S), .Y(
        early_flags_pmux_63_1_0_y0_8), .FCO(
        early_flags_pmux_63_1_0_co0_9));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[3]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[3]), .C(
        un10_early_flags[3]), .Y(late_flags_7_fast_Z[3]));
    SLE early_cur_set (.D(early_val_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_cur_set_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(early_cur_set_Z));
    SLE \retrain_reg[1]  (.D(retrain_reg_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(retrain_reg_Z[1]));
    CFG4 #( .INIT(16'h0020) )  bitalign_curr_state161 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state161_2_Z), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state161_Z));
    SLE \late_flags[99]  (.D(late_flags_7_fast_Z[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[99]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[6]  (.A(
        tapcnt_final_Z[6]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[6]), .Y(
        tapcnt_final_13_Z[6]));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_0_0 (.A(
        tapcnt_final_upd_Z[0]), .B(tapcnt_final_Z[0]), .C(tap_cnt_Z[0])
        , .D(N_1416), .Y(bitalign_curr_state61_0));
    CFG4 #( .INIT(16'h0001) )  calc_done25_177 (.A(early_flags_Z[51]), 
        .B(early_flags_Z[50]), .C(early_flags_Z[49]), .D(
        early_flags_Z[48]), .Y(calc_done25_177_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[88]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[88]), .C(
        un10_early_flags[88]), .Y(late_flags_7_fast_Z[88]));
    CFG2 #( .INIT(4'hE) )  un34lto7_3 (.A(un16_tapcnt_final_6), .B(
        un16_tapcnt_final_7), .Y(un34lto7_3_Z));
    SLE \rst_cnt[8]  (.D(rst_cnt_s[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[8]));
    CFG4 #( .INIT(16'h0053) )  \bitalign_curr_state_34_4_0_.m49  (.A(
        N_9), .B(N_11), .C(rx_err_Z), .D(bitalign_curr_state_Z[1]), .Y(
        N_50));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[4]), .D(
        late_flags_Z[68]), .FCI(late_flags_pmux_63_1_1_co1_4), .S(
        late_flags_pmux_63_1_1_wmux_11_S), .Y(
        late_flags_pmux_63_1_1_y0_4), .FCO(
        late_flags_pmux_63_1_1_co0_5));
    SLE \late_flags[103]  (.D(late_flags_7_fast_Z[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[103]));
    CFG4 #( .INIT(16'h0010) )  bitalign_curr_state148 (.A(
        bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state148_2_Z), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state148_Z));
    CFG3 #( .INIT(8'hF6) )  \wait_cnt_4[0]  (.A(
        bitalign_curr_state152_3_Z), .B(wait_cnt_Z[0]), .C(
        un1_restart_trng_fg_Z), .Y(wait_cnt_4_Z[0]));
    CFG2 #( .INIT(4'hD) )  bit_align_done_0_sqmuxa_3_i (.A(
        bit_align_done_0_sqmuxa_3_1_Z), .B(bit_align_done_0_sqmuxa_2_Z)
        , .Y(bit_align_done_0_sqmuxa_3_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[33]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[33]), .C(
        un10_early_flags[33]), .Y(early_flags_7_fast_Z[33]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[3]  (.A(
        tapcnt_final_Z[3]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[3]), .Y(
        tapcnt_final_13_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[51]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[51]), .C(
        un10_early_flags[51]), .Y(early_flags_7_fast_Z[51]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[16]), 
        .D(early_flags_Z[80]), .FCI(early_flags_pmux_63_1_1_co1), .S(
        early_flags_pmux_63_1_1_wmux_1_S), .Y(
        early_flags_pmux_63_1_1_y0_0), .FCO(
        early_flags_pmux_63_1_1_co0_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[94]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[94]), .C(
        un10_early_flags[94]), .Y(early_flags_7_fast_Z[94]));
    CFG4 #( .INIT(16'h3332) )  bit_align_start_RNO (.A(sig_re_train_Z), 
        .B(restart_trng_fg_i), .C(bit_align_done_0_sqmuxa_2_Z), .D(
        bitalign_curr_state_1_sqmuxa_4_Z), .Y(N_1439_i));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[90]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[90]), .C(
        un10_early_flags[90]), .Y(late_flags_7_fast_Z[90]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[35]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[35]), .C(
        un10_early_flags[35]), .Y(late_flags_7_fast_Z[35]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_122 (.A(tap_cnt_Z[2]), 
        .B(un10_early_flags_1_Z[10]), .C(un10_early_flags_1_Z[64]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[122]));
    CFG4 #( .INIT(16'h2772) )  \tapcnt_final_13_RNO_0[6]  (.A(
        tapcnt_final_3_sqmuxa_Z), .B(late_val_Z[6]), .C(
        un1_no_early_no_late_val_end1_1_1_Z[6]), .D(
        un1_no_early_no_late_val_st1_1_1[6]), .Y(
        tapcnt_final_13_m1_axb_6_1));
    SLE \early_flags[107]  (.D(early_flags_7_fast_Z[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[107]));
    CFG3 #( .INIT(8'h10) )  bitalign_curr_state_2_sqmuxa_4_0_0 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[1]), .C(
        bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state_2_sqmuxa_4_0_0_Z));
    CFG4 #( .INIT(16'h8000) )  reset_dly_fg4 (.A(rst_cnt_Z[0]), .B(
        reset_dly_fg4_8_Z), .C(rst_cnt_Z[1]), .D(reset_dly_fg4_4_Z), 
        .Y(reset_dly_fg4_Z));
    SLE \late_flags[101]  (.D(late_flags_7_fast_Z[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[101]));
    CFG1 #( .INIT(2'h1) )  tapcnt_final_upd_8_s_6_RNO (.A(
        mv_dn_fg_0_sqmuxa_i_o2_Z), .Y(N_12_i));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[25]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[25]), .C(
        un10_early_flags[25]), .Y(late_flags_7_fast_Z[25]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_3_0 (.A(
        emflag_cnt_Z[3]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[3]), .D(GND), .FCI(early_late_diff_8_cry_2), .S(
        early_late_diff_8[3]), .Y(early_late_diff_8_cry_3_0_Y), .FCO(
        early_late_diff_8_cry_3));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[2]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[2]), .C(
        un10_early_flags[2]), .Y(early_flags_7_fast_Z[2]));
    SLE \early_val[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[2]));
    CFG4 #( .INIT(16'hCECC) )  mv_dn_fg_0_sqmuxa_i_0 (.A(N_98), .B(
        mv_dn_fg_0_sqmuxa_i_o2_Z), .C(mv_dn_fg_Z), .D(mv_up_fg_Z), .Y(
        mv_dn_fg_0_sqmuxa_i_0_Z));
    SLE \no_early_no_late_val_st2[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[4]));
    SLE \tap_cnt[2]  (.D(N_28_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[2]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_162 (.A(early_flags_Z[127]), 
        .B(early_flags_Z[126]), .C(early_flags_Z[125]), .D(
        early_flags_Z[124]), .Y(calc_done25_162_Z));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_64_2_0 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[5]), .Y(
        un10_early_flags_2_0[64]));
    SLE bit_align_done (.D(bit_align_done_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        bit_align_done_0_sqmuxa_3_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(bit_align_done_Z)
        );
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[4]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[4]), .C(
        un10_early_flags[4]), .Y(late_flags_7_fast_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[3]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[3]), .C(
        un10_early_flags[3]), .Y(early_flags_7_fast_Z[3]));
    CFG3 #( .INIT(8'h73) )  no_early_no_late_val_st1_0_sqmuxa_i (.A(
        un1_early_flags_pmux_1_Z), .B(early_late_diff_0_sqmuxa_1_0_Z), 
        .C(emflag_cnt_0_sqmuxa), .Y(
        no_early_no_late_val_st1_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[41]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[41]), .C(
        un10_early_flags[41]), .Y(early_flags_7_fast_Z[41]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_175 (.A(early_flags_Z[75]), 
        .B(early_flags_Z[74]), .C(early_flags_Z[73]), .D(
        early_flags_Z[72]), .Y(calc_done25_175_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[102]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[102]), .C(
        un10_early_flags[102]), .Y(late_flags_7_fast_Z[102]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[11]), 
        .D(early_flags_Z[75]), .FCI(early_flags_pmux_126_1_0_co1_0), 
        .S(early_flags_pmux_126_1_0_wmux_3_S), .Y(
        early_flags_pmux_126_1_0_y0_1), .FCO(
        early_flags_pmux_126_1_0_co0_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[28]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[28]), .C(
        un10_early_flags[28]), .Y(early_flags_7_fast_Z[28]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_148 (.A(late_flags_Z[39]), 
        .B(late_flags_Z[38]), .C(late_flags_Z[37]), .D(
        late_flags_Z[36]), .Y(calc_done25_148_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[6]), .D(
        late_flags_Z[70]), .FCI(late_flags_pmux_63_1_0_co1_4), .S(
        late_flags_pmux_63_1_0_wmux_11_S), .Y(
        late_flags_pmux_63_1_0_y0_4), .FCO(
        late_flags_pmux_63_1_0_co0_5));
    CFG3 #( .INIT(8'hD0) )  early_flags_0_sqmuxa_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(BIT_ALGN_ERR_0_c), .C(
        bitalign_curr_state149_Z), .Y(early_flags_0_sqmuxa_1_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[88]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[88]), .C(
        un10_early_flags[88]), .Y(early_flags_7_fast_Z[88]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_0_wmux_20 (.A(
        late_flags_pmux_126_1_0_y0_8), .B(late_flags_pmux_126_1_0_y3_0)
        , .C(late_flags_pmux_126_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_0_co0_9), .S(
        late_flags_pmux_126_1_0_wmux_20_S), .Y(
        late_flags_pmux_126_1_0_0_y21), .FCO(
        late_flags_pmux_126_1_0_co1_9));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state148_4_1 (.A(
        bitalign_curr_state164_Z), .B(bitalign_curr_state162_Z), .C(
        bitalign_curr_state163_Z), .Y(un1_bitalign_curr_state148_4_1_Z)
        );
    CFG3 #( .INIT(8'hCE) )  mv_up_fg_0_sqmuxa_i_0 (.A(N_98), .B(
        mv_dn_fg_0_sqmuxa_i_o2_Z), .C(mv_up_fg_Z), .Y(
        mv_up_fg_0_sqmuxa_i_0_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[25]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[25]), .C(
        un10_early_flags[25]), .Y(early_flags_7_fast_Z[25]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[45]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[45]), .C(
        un10_early_flags[45]), .Y(late_flags_7_fast_Z[45]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[2]  (.A(
        tapcnt_final_Z[2]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[2]), .Y(
        tapcnt_final_13_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[85]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[85]), .C(
        un10_early_flags[85]), .Y(early_flags_7_fast_Z[85]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[30]), 
        .D(early_flags_Z[94]), .FCI(early_flags_pmux_63_1_0_co1_7), .S(
        early_flags_pmux_63_1_0_wmux_17_S), .Y(
        early_flags_pmux_63_1_0_y0_7), .FCO(
        early_flags_pmux_63_1_0_co0_8));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_0_wmux_8 (.A(
        early_flags_pmux_63_1_0_y0_3), .B(early_flags_pmux_63_1_0_0_y3)
        , .C(early_flags_pmux_63_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co0_3), .S(
        early_flags_pmux_63_1_0_wmux_8_S), .Y(
        early_flags_pmux_63_1_0_0_y9), .FCO(
        early_flags_pmux_63_1_0_co1_3));
    CFG3 #( .INIT(8'h08) )  bitalign_curr_state160 (.A(i22_mux_1), .B(
        bitalign_curr_state152_1_Z), .C(bitalign_curr_state_Z[4]), .Y(
        bitalign_curr_state160_Z));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_5 (.A(
        un10_tapcnt_final_5), .B(un16_tapcnt_final_5), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_4_Z), .S(
        un10_tapcnt_final_cry_5_S), .Y(un10_tapcnt_final_cry_5_Y), 
        .FCO(un10_tapcnt_final_cry_5_Z));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_6_2 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_2_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[68]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[68]), .C(
        un10_early_flags[68]), .Y(early_flags_7_fast_Z[68]));
    SLE \early_flags[89]  (.D(early_flags_7_fast_Z[89]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[89]));
    CFG2 #( .INIT(4'h1) )  \bitalign_curr_state_34_4_0_.m75  (.A(
        N_119_mux), .B(bitalign_curr_state_Z[0]), .Y(N_76_0));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_6 (.A(
        un16_tapcnt_final_6), .B(un10_tapcnt_final_6), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_5_Z), .S(
        un16_tapcnt_final_cry_6_S), .Y(un16_tapcnt_final_cry_6_Y), 
        .FCO(un16_tapcnt_final_cry_6_Z));
    CFG4 #( .INIT(16'h5554) )  tapcnt_final_1_sqmuxa_2_RNI2NBR (.A(
        restart_trng_fg_i), .B(tapcnt_final_1_sqmuxa_2_Z), .C(
        tapcnt_final_2_sqmuxa_Z), .D(tapcnt_final_3_sqmuxa_Z), .Y(
        un1_bitalign_curr_state169_12_sn));
    CFG4 #( .INIT(16'h0001) )  calc_done25_188 (.A(early_flags_Z[7]), 
        .B(early_flags_Z[6]), .C(early_flags_Z[5]), .D(
        early_flags_Z[4]), .Y(calc_done25_188_Z));
    CFG4 #( .INIT(16'hFFF8) )  un1_early_last_set_1_sqmuxa_1_1_tz (.A(
        bitalign_curr_state160_Z), .B(early_cur_set_Z), .C(
        emflag_cnt_0_sqmuxa), .D(bitalign_curr_state159_Z), .Y(
        un1_early_last_set_1_sqmuxa_1_1_tz_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[3]), .D(
        late_flags_Z[67]), .FCI(VCC), .S(
        late_flags_pmux_126_1_0_0_wmux_S), .Y(
        late_flags_pmux_126_1_0_0_y0), .FCO(
        late_flags_pmux_126_1_0_0_co0));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_2_0 (.A(
        emflag_cnt_Z[2]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[2]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_1), .S(
        noearly_nolate_diff_nxt_8[2]), .Y(
        noearly_nolate_diff_nxt_8_cry_2_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_2));
    SLE \noearly_nolate_diff_start[1]  (.D(
        noearly_nolate_diff_start_7[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_1));
    SLE \late_flags[50]  (.D(late_flags_RNO_Z[50]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[50]));
    CFG4 #( .INIT(16'h4073) )  \bitalign_curr_state_34_4_0_.m101  (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        N_100_0), .D(m101_1_1), .Y(N_102));
    CFG4 #( .INIT(16'h0001) )  calc_done25_166 (.A(early_flags_Z[111]), 
        .B(early_flags_Z[110]), .C(early_flags_Z[109]), .D(
        early_flags_Z[108]), .Y(calc_done25_166_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[65]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[65]), .C(
        un10_early_flags[65]), .Y(early_flags_7_fast_Z[65]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_47 (.A(
        un10_early_flags_47_0_Z), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[47]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_138 (.A(late_flags_Z[95]), 
        .B(late_flags_Z[94]), .C(late_flags_Z[93]), .D(
        late_flags_Z[92]), .Y(calc_done25_138_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[52]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[52]), .C(
        un10_early_flags[52]), .Y(late_flags_7_fast_Z[52]));
    CFG4 #( .INIT(16'h8000) )  early_flags_dec_127_4 (.A(
        emflag_cnt_Z[4]), .B(emflag_cnt_Z[3]), .C(emflag_cnt_Z[6]), .D(
        emflag_cnt_Z[5]), .Y(early_flags_dec_127_4_Z));
    CFG4 #( .INIT(16'h8000) )  reset_dly_fg4_8 (.A(rst_cnt_Z[9]), .B(
        rst_cnt_Z[7]), .C(rst_cnt_Z[6]), .D(reset_dly_fg4_6_Z), .Y(
        reset_dly_fg4_8_Z));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNICU2D1[3]  (.A(early_val_Z[3])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[3]), .Y(
        early_val_RNICU2D1_Z[3]));
    CFG3 #( .INIT(8'hEC) )  rx_trng_done1_1_sqmuxa_i_o2 (.A(
        un1_rx_BIT_ALGN_START), .B(bitalign_curr_state12_Z), .C(
        un1_retrain_adj_tap_i), .Y(N_61));
    CFG2 #( .INIT(4'h7) )  \bitalign_curr_state_34_4_0_.N_29_i  (.A(
        bitalign_curr_state41_Z), .B(bitalign_curr_state_Z[0]), .Y(
        N_29_i));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_33 (.A(tap_cnt_Z[0]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_2_0[32]), .Y(un10_early_flags[33]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[120]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[120]), .C(
        un10_early_flags[120]), .Y(early_flags_7_fast_Z[120]));
    SLE \late_flags[126]  (.D(late_flags_7_fast_Z[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[126]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[70]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[70]), .C(
        un10_early_flags[70]), .Y(early_flags_7_fast_Z[70]));
    SLE \early_flags[28]  (.D(early_flags_7_fast_Z[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[28]));
    SLE \restart_edge_reg[1]  (.D(restart_edge_reg_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[1]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_63_1_0_wmux_8 (.A(
        late_flags_pmux_63_1_0_y0_3), .B(late_flags_pmux_63_1_0_0_y3), 
        .C(late_flags_pmux_63_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co0_3), .S(
        late_flags_pmux_63_1_0_wmux_8_S), .Y(
        late_flags_pmux_63_1_0_0_y9), .FCO(
        late_flags_pmux_63_1_0_co1_3));
    SLE \early_late_diff[7]  (.D(early_late_diff_8[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[7]));
    SLE \no_early_no_late_val_st1[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[5]));
    SLE \early_flags[44]  (.D(early_flags_7_fast_Z[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[44]));
    SLE \early_flags[121]  (.D(early_flags_7_fast_Z[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[121]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNI8CA5K[5]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIROIR_Z[5]), .B(
        early_val_RNII43D1_Z[5]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[5]), .FCI(tapcnt_final_13_m1_cry_4), .S(
        tapcnt_final_13_m1[5]), .Y(early_val_RNI8CA5K_Y[5]), .FCO(
        tapcnt_final_13_m1_cry_5));
    CFG3 #( .INIT(8'hE4) )  \late_flags_RNO[50]  (.A(N_209), .B(
        EYE_MONITOR_LATE_net_0_0), .C(late_flags_Z[50]), .Y(
        late_flags_RNO_Z[50]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[29]), 
        .D(early_flags_Z[93]), .FCI(early_flags_pmux_126_1_1_co1_7), 
        .S(early_flags_pmux_126_1_1_wmux_17_S), .Y(
        early_flags_pmux_126_1_1_y0_7), .FCO(
        early_flags_pmux_126_1_1_co0_8));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_127_1_0_wmux_0 (.A(
        late_flags_pmux_127_1_0_y0), .B(emflag_cnt_Z[0]), .C(
        late_flags_pmux_126_1_1_wmux_10_Y), .D(
        late_flags_pmux_126_1_0_wmux_10_Y), .FCI(
        late_flags_pmux_127_1_0_co0), .S(
        late_flags_pmux_127_1_0_wmux_0_S), .Y(late_flags_pmux), .FCO(
        late_flags_pmux_127_1_0_co1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[37]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[37]), .C(
        un10_early_flags[37]), .Y(late_flags_7_fast_Z[37]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_54 (.A(tap_cnt_Z[6]), 
        .B(un10_early_flags_2_Z[6]), .C(un10_early_flags_1_Z[6]), .D(
        un10_early_flags_1_Z[48]), .Y(un10_early_flags[54]));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[2]  (.A(N_78), .B(N_63_0), .Y(
        N_28_i));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_7 (.A(
        un10_tapcnt_final_7), .B(early_late_diff_Z[7]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_6_Z), .S(
        un1_early_late_diff_cry_7_S), .Y(un1_early_late_diff_cry_7_Y), 
        .FCO(un1_early_late_diff_cry_7_Z));
    CFG3 #( .INIT(8'hFB) )  \tap_cnt_17_i_o2_0[6]  (.A(
        un1_early_flags_1_sqmuxa_i), .B(
        bitalign_curr_state_0_sqmuxa_10), .C(
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), .Y(N_60));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[22]), 
        .D(late_flags_Z[86]), .FCI(late_flags_pmux_63_1_0_co1_5), .S(
        late_flags_pmux_63_1_0_wmux_13_S), .Y(
        late_flags_pmux_63_1_0_y0_5), .FCO(
        late_flags_pmux_63_1_0_co0_6));
    SLE \early_flags[99]  (.D(early_flags_7_fast_Z[99]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[99]));
    CFG2 #( .INIT(4'h2) )  rx_trng_done_1_sqmuxa (.A(
        bitalign_curr_state164_Z), .B(bitalign_curr_state41_Z), .Y(
        rx_trng_done_1_sqmuxa_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[1]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[1]), .C(
        un10_early_flags[1]), .Y(early_flags_7_fast_Z[1]));
    SLE \early_flags[100]  (.D(early_flags_7_fast_Z[100]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[100]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_0 (.A(
        un16_tapcnt_final_0), .B(early_late_diff_Z[0]), .C(GND), .D(
        GND), .FCI(GND), .S(un1_early_late_diff_1_cry_0_S), .Y(
        un1_early_late_diff_1_cry_0_Y), .FCO(
        un1_early_late_diff_1_cry_0_Z));
    SLE \timeout_cnt[5]  (.D(timeout_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(timeout_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(timeout_cnt_Z[5]));
    SLE \emflag_cnt[1]  (.D(emflag_cnt_s[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[1]));
    SLE \early_flags[123]  (.D(early_flags_7_fast_Z[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[123]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[98]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[98]), .C(
        un10_early_flags[98]), .Y(late_flags_7_fast_Z[98]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[27]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[27]), .C(
        un10_early_flags[27]), .Y(late_flags_7_fast_Z[27]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[6]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[6]), .C(
        un10_early_flags[6]), .Y(late_flags_7_fast_Z[6]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_18 (.A(
        early_flags_pmux_126_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[61]), .D(early_flags_Z[125]), .FCI(
        early_flags_pmux_126_1_1_co0_8), .S(
        early_flags_pmux_126_1_1_wmux_18_S), .Y(
        early_flags_pmux_126_1_1_y7_0), .FCO(
        early_flags_pmux_126_1_1_co1_8));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_23 (.A(
        un10_early_flags_2_0[16]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[20]), .Y(un10_early_flags[23]));
    SLE \late_flags[27]  (.D(late_flags_7_fast_Z[27]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[27]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[2]), .D(
        late_flags_Z[66]), .FCI(VCC), .S(
        late_flags_pmux_63_1_0_0_wmux_S), .Y(
        late_flags_pmux_63_1_0_0_y0), .FCO(
        late_flags_pmux_63_1_0_0_co0));
    SLE \late_flags[60]  (.D(late_flags_7_fast_Z[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[60]));
    CFG2 #( .INIT(4'hE) )  un1_bitalign_curr_state_13_1 (.A(
        early_flags_0_sqmuxa_1_Z), .B(bitalign_curr_state_Z[4]), .Y(
        un1_bitalign_curr_state_13_1_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_142 (.A(late_flags_Z[79]), 
        .B(late_flags_Z[78]), .C(late_flags_Z[77]), .D(
        late_flags_Z[76]), .Y(calc_done25_142_Z));
    CFG2 #( .INIT(4'h9) )  un1_bitalign_curr_state151 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state151_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_64 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_2_0[64]), .C(
        un10_early_flags_2_Z[8]), .Y(un10_early_flags[64]));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_0_wmux_8 (.A(
        early_flags_pmux_126_1_0_y0_3), .B(
        early_flags_pmux_126_1_0_0_y3), .C(
        early_flags_pmux_126_1_0_0_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_0_co0_3), .S(
        early_flags_pmux_126_1_0_wmux_8_S), .Y(
        early_flags_pmux_126_1_0_0_y9), .FCO(
        early_flags_pmux_126_1_0_co1_3));
    CFG2 #( .INIT(4'h8) )  calc_done25_209 (.A(calc_done25_162_Z), .B(
        calc_done25_163_Z), .Y(calc_done25_209_Z));
    SLE \early_flags[2]  (.D(early_flags_7_fast_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[2]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_46 (.A(
        un10_early_flags_3_Z[46]), .B(tap_cnt_Z[6]), .C(
        un10_early_flags_1_Z[6]), .D(un10_early_flags_1_Z[40]), .Y(
        un10_early_flags[46]));
    SLE \late_flags[107]  (.D(late_flags_7_fast_Z[107]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[107]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[122]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[122]), .C(
        un10_early_flags[122]), .Y(late_flags_7_fast_Z[122]));
    SLE \early_flags[46]  (.D(early_flags_7_fast_Z[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[46]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_235 (.A(calc_done25_175_Z), 
        .B(calc_done25_174_Z), .C(calc_done25_173_Z), .D(
        calc_done25_172_Z), .Y(calc_done25_235_Z));
    SLE \early_flags[47]  (.D(early_flags_7_fast_Z[47]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[47]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[72]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[72]), .C(
        un10_early_flags[72]), .Y(late_flags_7_fast_Z[72]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[118]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[118]), .C(
        un10_early_flags[118]), .Y(late_flags_7_fast_Z[118]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_9 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_63_1_1_co1_3), .S(
        late_flags_pmux_63_1_1_wmux_9_S), .Y(
        late_flags_pmux_63_1_1_wmux_9_Y), .FCO(
        late_flags_pmux_63_1_1_co0_4));
    SLE \late_flags[77]  (.D(late_flags_7_fast_Z[77]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[77]));
    SLE \early_late_diff[5]  (.D(early_late_diff_8[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[74]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[74]), .C(
        un10_early_flags[74]), .Y(early_flags_7_fast_Z[74]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_182 (.A(early_flags_Z[47]), 
        .B(early_flags_Z[46]), .C(early_flags_Z[45]), .D(
        early_flags_Z[44]), .Y(calc_done25_182_Z));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_7 (.A(
        late_flags_pmux_126_1_1_y7), .B(late_flags_pmux_126_1_1_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co1_2), .S(
        late_flags_pmux_126_1_1_wmux_7_S), .Y(
        late_flags_pmux_126_1_1_y0_3), .FCO(
        late_flags_pmux_126_1_1_co0_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[47]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[47]), .C(
        un10_early_flags[47]), .Y(late_flags_7_fast_Z[47]));
    SLE \early_flags[41]  (.D(early_flags_7_fast_Z[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[41]));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_114 (.A(tap_cnt_Z[3]), 
        .B(N_1499), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[114]));
    CFG4 #( .INIT(16'h8000) )  rx_BIT_ALGN_ERR (.A(timeout_cnt_Z[4]), 
        .B(timeout_cnt_Z[5]), .C(rx_BIT_ALGN_ERR_4_Z), .D(
        rx_BIT_ALGN_ERR_3_Z), .Y(BIT_ALGN_ERR_0_c));
    CFG4 #( .INIT(16'h0001) )  calc_done25_132 (.A(late_flags_Z[103]), 
        .B(late_flags_Z[102]), .C(late_flags_Z[101]), .D(
        late_flags_Z[100]), .Y(calc_done25_132_Z));
    CFG2 #( .INIT(4'hE) )  un1_restart_trng_fg_10_0 (.A(
        un1_restart_trng_fg_10_sn_1), .B(tap_cnt_0_sqmuxa_1_Z), .Y(
        un1_restart_trng_fg_10_0_Z));
    CFG4 #( .INIT(16'hBFFF) )  \late_flags_7_i_o4[50]  (.A(
        tap_cnt_Z[0]), .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[48]), 
        .D(un10_early_flags_1_Z[48]), .Y(N_209));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_72 (.A(
        un10_early_flags_2_0[72]), .B(un10_early_flags_1_Z[0]), .C(
        un10_early_flags_1_Z[72]), .Y(un10_early_flags[72]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_16 (.A(
        early_flags_pmux_63_1_1_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[44]), .D(early_flags_Z[108]), .FCI(
        early_flags_pmux_63_1_1_co0_7), .S(
        early_flags_pmux_63_1_1_wmux_16_S), .Y(
        early_flags_pmux_63_1_1_y5_0), .FCO(
        early_flags_pmux_63_1_1_co1_7));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_14 (.A(
        early_flags_pmux_63_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[52]), .D(early_flags_Z[116]), .FCI(
        early_flags_pmux_63_1_1_co0_6), .S(
        early_flags_pmux_63_1_1_wmux_14_S), .Y(
        early_flags_pmux_63_1_1_y3_0), .FCO(
        early_flags_pmux_63_1_1_co1_6));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[3]), 
        .D(early_flags_Z[67]), .FCI(VCC), .S(
        early_flags_pmux_126_1_0_0_wmux_S), .Y(
        early_flags_pmux_126_1_0_0_y0), .FCO(
        early_flags_pmux_126_1_0_0_co0));
    SLE \late_flags[86]  (.D(late_flags_7_fast_Z[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[86]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_146 (.A(late_flags_Z[51]), 
        .B(late_flags_Z[50]), .C(late_flags_Z[49]), .D(
        late_flags_Z[48]), .Y(calc_done25_146_Z));
    SLE \noearly_nolate_diff_nxt[5]  (.D(noearly_nolate_diff_nxt_8[5]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_5));
    SLE \early_late_diff[2]  (.D(early_late_diff_8[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[2]));
    SLE \late_flags[37]  (.D(late_flags_7_fast_Z[37]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[37]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[23]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[23]), .C(
        un10_early_flags[23]), .Y(early_flags_7_fast_Z[23]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_6 (.A(
        late_flags_pmux_63_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[56]), .D(late_flags_Z[120]), .FCI(
        late_flags_pmux_63_1_1_co0_2), .S(
        late_flags_pmux_63_1_1_wmux_6_S), .Y(late_flags_pmux_63_1_1_y7)
        , .FCO(late_flags_pmux_63_1_1_co1_2));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[83]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[83]), .C(
        un10_early_flags[83]), .Y(early_flags_7_fast_Z[83]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNI9AK2A[2]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNILIIR_Z[2]), .B(
        early_val_RNI9R2D1_Z[2]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[2]), .FCI(tapcnt_final_13_m1_cry_1), .S(
        tapcnt_final_13_m1[2]), .Y(early_val_RNI9AK2A_Y[2]), .FCO(
        tapcnt_final_13_m1_cry_2));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_4 (.A(
        un10_tapcnt_final_4), .B(early_late_diff_Z[4]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_3_Z), .S(
        un1_early_late_diff_cry_4_S), .Y(un1_early_late_diff_cry_4_Y), 
        .FCO(un1_early_late_diff_cry_4_Z));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_4_0 (.A(
        emflag_cnt_Z[4]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[4]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_3), .S(
        noearly_nolate_diff_nxt_8[4]), .Y(
        noearly_nolate_diff_nxt_8_cry_4_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_4));
    CFG3 #( .INIT(8'h80) )  rx_BIT_ALGN_LOAD_0_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(tap_cnt_0_sqmuxa_2_0), .C(
        un1_bitalign_curr_state152_Z), .Y(rx_BIT_ALGN_LOAD_0_sqmuxa_Z));
    SLE rx_BIT_ALGN_MOVE (.D(rx_BIT_ALGN_MOVE_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE));
    SLE \late_flags[16]  (.D(late_flags_7_fast_Z[16]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[16]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[12]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[12]), .C(
        un10_early_flags[12]), .Y(early_flags_7_fast_Z[12]));
    CFG4 #( .INIT(16'hAAEA) )  un1_restart_trng_fg (.A(
        restart_trng_fg_i), .B(bitalign_curr_state148_2_Z), .C(
        bitalign_curr_state_Z[1]), .D(bitalign_curr_state_Z[0]), .Y(
        un1_restart_trng_fg_Z));
    CFG4 #( .INIT(16'h8880) )  un1_early_late_diff_valid (.A(
        late_last_set_Z), .B(early_last_set_Z), .C(
        un2_early_late_diff_validlto7_2_Z), .D(
        un2_early_late_diff_validlt7), .Y(un1_early_late_diff_valid_Z));
    CFG4 #( .INIT(16'hFF13) )  un1_restart_trng_fg_6 (.A(
        bitalign_curr_state155_Z), .B(tapcnt_final_upd_2_sqmuxa), .C(
        mv_dn_fg_Z), .D(restart_trng_fg_i), .Y(un1_restart_trng_fg_6_Z)
        );
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[104]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[104]), .C(
        un10_early_flags[104]), .Y(late_flags_7_fast_Z[104]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[5]), 
        .D(early_flags_Z[69]), .FCI(early_flags_pmux_126_1_1_co1_4), 
        .S(early_flags_pmux_126_1_1_wmux_11_S), .Y(
        early_flags_pmux_126_1_1_y0_4), .FCO(
        early_flags_pmux_126_1_1_co0_5));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[63]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[63]), .C(
        un10_early_flags[63]), .Y(early_flags_7_fast_Z[63]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_186 (.A(early_flags_Z[31]), 
        .B(early_flags_Z[30]), .C(early_flags_Z[29]), .D(
        early_flags_Z[28]), .Y(calc_done25_186_Z));
    SLE \early_flags[30]  (.D(early_flags_7_fast_Z[30]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[30]));
    CFG3 #( .INIT(8'h08) )  mv_dn_fg_0_sqmuxa_i_a2_0 (.A(
        retrain_reg_Z[2]), .B(bitalign_curr_state148_Z), .C(
        BIT_ALGN_ERR_0_c), .Y(N_98));
    SLE \late_flags[55]  (.D(late_flags_7_fast_Z[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[55]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[6]  (.A(VCC), .B(
        rst_cnt_Z[6]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[5]), .S(
        rst_cnt_s[6]), .Y(rst_cnt_cry_Y_0[6]), .FCO(rst_cnt_cry_Z[6]));
    CFG2 #( .INIT(4'h4) )  reset_dly_fg4_4 (.A(reset_dly_fg_Z), .B(
        rst_cnt_Z[8]), .Y(reset_dly_fg4_4_Z));
    SLE \early_flags[55]  (.D(early_flags_7_fast_Z[55]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[55]));
    CFG4 #( .INIT(16'h353F) )  \bitalign_curr_state_34_4_0_.m50_1_1  (
        .A(bitalign_curr_state41_Z), .B(N_50), .C(
        bitalign_curr_state_Z[2]), .D(bitalign_curr_state_Z[0]), .Y(
        m50_1_1));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_4 (.A(
        early_flags_pmux_63_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[42]), .D(early_flags_Z[106]), .FCI(
        early_flags_pmux_63_1_0_co0_1), .S(
        early_flags_pmux_63_1_0_wmux_4_S), .Y(
        early_flags_pmux_63_1_0_0_y5), .FCO(
        early_flags_pmux_63_1_0_co1_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[98]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[98]), .C(
        un10_early_flags[98]), .Y(early_flags_7_fast_Z[98]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_136 (.A(late_flags_Z[87]), 
        .B(late_flags_Z[86]), .C(late_flags_Z[85]), .D(
        late_flags_Z[84]), .Y(calc_done25_136_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[54]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[54]), .C(
        un10_early_flags[54]), .Y(late_flags_7_fast_Z[54]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_104 (.A(
        un10_early_flags_1_Z[40]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[64]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[104]));
    SLE \tapcnt_final_upd[4]  (.D(tapcnt_final_upd_8[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[4]));
    SLE \late_flags[46]  (.D(late_flags_7_fast_Z[46]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[46]));
    ARI1 #( .INIT(20'h45500) )  early_late_diff_8_cry_0_0_cy (.A(VCC), 
        .B(un1_restart_trng_fg_5_Z), .C(GND), .D(GND), .FCI(VCC), .S(
        early_late_diff_8_cry_0_0_cy_S), .Y(
        early_late_diff_8_cry_0_0_cy_Y), .FCO(
        early_late_diff_8_cry_0_0_cy_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[95]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[95]), .C(
        un10_early_flags[95]), .Y(early_flags_7_fast_Z[95]));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_1_wmux_20 (.A(
        late_flags_pmux_126_1_1_y0_8), .B(late_flags_pmux_126_1_1_y3_0)
        , .C(late_flags_pmux_126_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co0_9), .S(
        late_flags_pmux_126_1_1_wmux_20_S), .Y(
        late_flags_pmux_126_1_1_y21), .FCO(
        late_flags_pmux_126_1_1_co1_9));
    CFG2 #( .INIT(4'h1) )  early_late_diff_0_sqmuxa_1_0 (.A(
        un1_tap_cnt_0_sqmuxa_6_0), .B(restart_trng_fg_i), .Y(
        early_late_diff_0_sqmuxa_1_0_Z));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_0 (.A(
        early_flags_pmux_126_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[35]), .D(early_flags_Z[99]), .FCI(
        early_flags_pmux_126_1_0_0_co0), .S(
        early_flags_pmux_126_1_0_wmux_0_S), .Y(
        early_flags_pmux_126_1_0_0_y1), .FCO(
        early_flags_pmux_126_1_0_0_co1));
    SLE \restart_edge_reg[3]  (.D(restart_edge_reg_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[3]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_14 (.A(
        late_flags_pmux_126_1_0_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[55]), .D(late_flags_Z[119]), .FCI(
        late_flags_pmux_126_1_0_co0_6), .S(
        late_flags_pmux_126_1_0_wmux_14_S), .Y(
        late_flags_pmux_126_1_0_y3_0), .FCO(
        late_flags_pmux_126_1_0_co1_6));
    CFG2 #( .INIT(4'hE) )  un1_early_flags_pmux_1 (.A(early_flags_pmux)
        , .B(late_flags_pmux), .Y(un1_early_flags_pmux_1_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_18 (.A(
        late_flags_pmux_126_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[61]), .D(late_flags_Z[125]), .FCI(
        late_flags_pmux_126_1_1_co0_8), .S(
        late_flags_pmux_126_1_1_wmux_18_S), .Y(
        late_flags_pmux_126_1_1_y7_0), .FCO(
        late_flags_pmux_126_1_1_co1_8));
    SLE \emflag_cnt[0]  (.D(emflag_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_18 (.A(
        late_flags_pmux_63_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[60]), .D(late_flags_Z[124]), .FCI(
        late_flags_pmux_63_1_1_co0_8), .S(
        late_flags_pmux_63_1_1_wmux_18_S), .Y(
        late_flags_pmux_63_1_1_y7_0), .FCO(
        late_flags_pmux_63_1_1_co1_8));
    SLE \noearly_nolate_diff_start[3]  (.D(
        noearly_nolate_diff_start_7[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_3));
    SLE \late_flags[81]  (.D(late_flags_7_fast_Z[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[81]));
    CFG4 #( .INIT(16'hCCEF) )  \emflag_cnt_cry_cy_RNO[0]  (.A(
        bitalign_curr_state_Z[0]), .B(restart_trng_fg_i), .C(
        bitalign_curr_state_Z[4]), .D(bitalign_curr_state_Z[2]), .Y(
        un1_restart_trng_fg_9_0_443_0));
    CFG4 #( .INIT(16'hAABA) )  rx_trng_done1_0_sqmuxa_i (.A(
        restart_trng_fg_i), .B(un1_bitalign_curr_state_16_1_Z), .C(
        N_52), .D(early_flags_0_sqmuxa_1_Z), .Y(
        rx_trng_done1_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[30]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[30]), .C(
        un10_early_flags[30]), .Y(late_flags_7_fast_Z[30]));
    SLE \early_flags[60]  (.D(early_flags_7_fast_Z[60]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[60]));
    ARI1 #( .INIT(20'h0F588) )  
        \bitalign_curr_state_34_4_0_.m74_2_1_1_wmux_0  (.A(
        m74_2_1_1_1_y0), .B(bitalign_curr_state_Z[1]), .C(N_29_i), .D(
        N_116_mux), .FCI(m74_2_1_1_1_co0), .S(m74_2_1_1_wmux_0_S), .Y(
        N_75_0), .FCO(m74_2_1_1_1_co1));
    CFG4 #( .INIT(16'h0001) )  calc_done25_164 (.A(early_flags_Z[103]), 
        .B(early_flags_Z[102]), .C(early_flags_Z[101]), .D(
        early_flags_Z[100]), .Y(calc_done25_164_Z));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_57 (.A(
        un10_early_flags_1_Z[9]), .B(tap_cnt_Z[6]), .C(
        un10_early_flags_1_Z[48]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[57]));
    CFG3 #( .INIT(8'h08) )  \bitalign_curr_state_34_4_0_.m110  (.A(
        bitalign_curr_state161_2_Z), .B(N_76_0), .C(
        bitalign_curr_state_Z[3]), .Y(N_130_mux));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_6 (.A(
        early_flags_pmux_126_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[59]), .D(early_flags_Z[123]), .FCI(
        early_flags_pmux_126_1_0_co0_2), .S(
        early_flags_pmux_126_1_0_wmux_6_S), .Y(
        early_flags_pmux_126_1_0_0_y7), .FCO(
        early_flags_pmux_126_1_0_co1_2));
    CFG4 #( .INIT(16'h0800) )  bitalign_curr_state_2_sqmuxa_4_0 (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .C(
        early_flags_dec[127]), .D(bitalign_curr_state_2_sqmuxa_4_0_0_Z)
        , .Y(emflag_cnt_0_sqmuxa));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[0]  (.A(
        no_early_no_late_val_end1_Z[0]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[0]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[0]));
    SLE \no_early_no_late_val_end2[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[0]));
    SLE \late_flags[65]  (.D(late_flags_7_fast_Z[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[65]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[20]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[20]), .C(
        un10_early_flags[20]), .Y(late_flags_7_fast_Z[20]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[116]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[116]), .C(
        un10_early_flags[116]), .Y(late_flags_7_fast_Z[116]));
    CFG3 #( .INIT(8'hFB) )  early_cur_set_0_sqmuxa_i (.A(
        un1_tap_cnt_0_sqmuxa_6_0), .B(early_cur_set_0_sqmuxa_1_Z), .C(
        early_val_0_sqmuxa_1_0_Z), .Y(early_cur_set_0_sqmuxa_i_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_112 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_1_Z[48]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[112]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[29]), 
        .D(late_flags_Z[93]), .FCI(late_flags_pmux_126_1_1_co1_7), .S(
        late_flags_pmux_126_1_1_wmux_17_S), .Y(
        late_flags_pmux_126_1_1_y0_7), .FCO(
        late_flags_pmux_126_1_1_co0_8));
    CFG4 #( .INIT(16'h0001) )  calc_done25_151 (.A(late_flags_Z[43]), 
        .B(late_flags_Z[42]), .C(late_flags_Z[41]), .D(
        late_flags_Z[40]), .Y(calc_done25_151_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[25]), 
        .D(early_flags_Z[89]), .FCI(early_flags_pmux_126_1_1_co1_1), 
        .S(early_flags_pmux_126_1_1_wmux_5_S), .Y(
        early_flags_pmux_126_1_1_y0_2), .FCO(
        early_flags_pmux_126_1_1_co0_2));
    CFG2 #( .INIT(4'h8) )  rx_BIT_ALGN_ERR_3 (.A(timeout_cnt_Z[6]), .B(
        timeout_cnt_Z[7]), .Y(rx_BIT_ALGN_ERR_3_Z));
    SLE \late_flags[11]  (.D(late_flags_7_fast_Z[11]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[11]));
    SLE \early_flags[32]  (.D(early_flags_7_fast_Z[32]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[32]));
    SLE \early_flags[7]  (.D(early_flags_7_fast_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[7]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_19 (.A(
        late_flags_pmux_63_1_0_y7_0), .B(late_flags_pmux_63_1_0_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_0_co1_8), .S(
        late_flags_pmux_63_1_0_wmux_19_S), .Y(
        late_flags_pmux_63_1_0_y0_8), .FCO(
        late_flags_pmux_63_1_0_co0_9));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[11]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[11]), .C(
        un10_early_flags[11]), .Y(late_flags_7_fast_Z[11]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_67 (.A(
        un10_early_flags_2_0[64]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_2_Z[67]), .Y(un10_early_flags[67]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[1]), 
        .D(early_flags_Z[65]), .FCI(VCC), .S(
        early_flags_pmux_126_1_1_wmux_S), .Y(
        early_flags_pmux_126_1_1_y0), .FCO(
        early_flags_pmux_126_1_1_co0));
    CFG4 #( .INIT(16'hAE00) )  tapcnt_final_2_sqmuxa (.A(calc_done28_Z)
        , .B(calc_done27_Z), .C(un10_tapcnt_final_cry_7_Z), .D(
        bitalign_curr_state162_Z), .Y(tapcnt_final_2_sqmuxa_Z));
    SLE \rst_cnt[7]  (.D(rst_cnt_s[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[7]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[103]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[103]), .C(
        un10_early_flags[103]), .Y(late_flags_7_fast_Z[103]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[6]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[6]), .C(
        un10_early_flags[6]), .Y(early_flags_7_fast_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[12]), 
        .D(early_flags_Z[76]), .FCI(early_flags_pmux_63_1_1_co1_6), .S(
        early_flags_pmux_63_1_1_wmux_15_S), .Y(
        early_flags_pmux_63_1_1_y0_6), .FCO(
        early_flags_pmux_63_1_1_co0_7));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIHEIR[0]  (.A(
        late_val_Z[0]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[0]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIHEIR_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[74]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[74]), .C(
        un10_early_flags[74]), .Y(late_flags_7_fast_Z[74]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[24]), 
        .D(late_flags_Z[88]), .FCI(late_flags_pmux_63_1_1_co1_1), .S(
        late_flags_pmux_63_1_1_wmux_5_S), .Y(
        late_flags_pmux_63_1_1_y0_2), .FCO(
        late_flags_pmux_63_1_1_co0_2));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_75 (.A(
        un10_early_flags_2_0[72]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[72]), .Y(un10_early_flags[75]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_121 (.A(
        un10_early_flags_1_Z[9]), .B(tap_cnt_Z[2]), .C(
        un10_early_flags_1_Z[48]), .D(un10_early_flags_2_Z[69]), .Y(
        un10_early_flags[121]));
    SLE \late_flags[41]  (.D(late_flags_7_fast_Z[41]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[41]));
    SLE \early_flags[125]  (.D(early_flags_7_fast_Z[125]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[125]));
    SLE \early_flags[48]  (.D(early_flags_7_fast_Z[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[48]));
    SLE \late_flags[23]  (.D(late_flags_7_fast_Z[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[23]));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_3_sqmuxa (.A(
        early_flags_1_sqmuxa_1_Z), .B(un1_rx_BIT_ALGN_START), .Y(
        tapcnt_final_upd_3_sqmuxa_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_99 (.A(
        un10_early_flags_1_Z[3]), .B(un10_early_flags_2_0[96]), .C(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[99]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_4_0 (.A(
        emflag_cnt_Z[4]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[4]), .D(GND), .FCI(early_late_diff_8_cry_3), .S(
        early_late_diff_8[4]), .Y(early_late_diff_8_cry_4_0_Y), .FCO(
        early_late_diff_8_cry_4));
    CFG4 #( .INIT(16'h8000) )  calc_done25_224 (.A(calc_done25_131_Z), 
        .B(calc_done25_130_Z), .C(calc_done25_129_Z), .D(
        calc_done25_128_Z), .Y(calc_done25_224_Z));
    SLE \late_flags[96]  (.D(late_flags_7_fast_Z[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[96]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[40]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[40]), .C(
        un10_early_flags[40]), .Y(late_flags_7_fast_Z[40]));
    CFG2 #( .INIT(4'h2) )  bitalign_curr_state_0_sqmuxa_10_0_a2 (.A(
        N_100), .B(un1_retrain_adj_tap_i), .Y(
        bitalign_curr_state_0_sqmuxa_10));
    SLE \early_flags[70]  (.D(early_flags_7_fast_Z[70]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[70]));
    SLE \early_flags[62]  (.D(early_flags_7_fast_Z[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[62]));
    SLE \early_flags[117]  (.D(early_flags_7_fast_Z[117]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[117]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_56 (.A(
        un10_early_flags_1_Z[32]), .B(tap_cnt_Z[6]), .C(
        un10_early_flags_1_Z[24]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[56]));
    SLE early_last_set (.D(early_last_set_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_last_set_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(early_last_set_Z)
        );
    CFG3 #( .INIT(8'hAB) )  tapcnt_final_upd_0_sqmuxa_i (.A(
        restart_trng_fg_i), .B(un1_bitalign_curr_state_13_1_Z), .C(
        un1_bitalign_curr_state_14_1_Z), .Y(
        tapcnt_final_upd_0_sqmuxa_i_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[124]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[124]), .C(
        un10_early_flags[124]), .Y(late_flags_7_fast_Z[124]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_0_0 (.A(
        emflag_cnt_Z[0]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[0]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_0_0_cy_Z), .S(
        noearly_nolate_diff_nxt_8[0]), .Y(
        noearly_nolate_diff_nxt_8_cry_0_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_0));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_126_1_0_wmux_20 (.A(
        early_flags_pmux_126_1_0_y0_8), .B(
        early_flags_pmux_126_1_0_y3_0), .C(
        early_flags_pmux_126_1_0_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_0_co0_9), .S(
        early_flags_pmux_126_1_0_wmux_20_S), .Y(
        early_flags_pmux_126_1_0_0_y21), .FCO(
        early_flags_pmux_126_1_0_co1_9));
    CFG4 #( .INIT(16'hFFFE) )  un1_bitalign_curr_state_15_3 (.A(
        rx_BIT_ALGN_DIR_1_sqmuxa_Z), .B(early_flags_0_sqmuxa_1_Z), .C(
        un1_bitalign_curr_state_15_0_Z), .D(early_flags_0_sqmuxa_Z), 
        .Y(un1_bitalign_curr_state_15_3_Z));
    CFG2 #( .INIT(4'h7) )  un10_early_flags_17_1_i (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[0]), .Y(N_1498));
    CFG4 #( .INIT(16'hA5EC) )  \tapcnt_final_13_1[0]  (.A(
        tapcnt_final_13_1_1_0_Z[0]), .B(tapcnt_final_13_Z[1]), .C(
        tapcnt_final_13_m0s2_Z), .D(un1_tapcnt_final_0_sqmuxa_Z), .Y(
        tapcnt_final_13_1_Z[0]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_102 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[96]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_2_Z[6]), .Y(
        un10_early_flags[102]));
    SLE rx_err (.D(N_1392), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        rx_err_0_sqmuxa_1_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC)
        , .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_err_Z));
    SLE \early_flags[85]  (.D(early_flags_7_fast_Z[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[85]));
    CFG4 #( .INIT(16'hFFFE) )  un34lto7 (.A(un16_tapcnt_final_4), .B(
        un16_tapcnt_final_5), .C(un34lto7_4_Z), .D(un34lto7_3_Z), .Y(
        un34));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[65]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[65]), .C(
        un10_early_flags[65]), .Y(late_flags_7_fast_Z[65]));
    CFG1 #( .INIT(2'h1) )  \cnt_RNO[0]  (.A(CO0_0), .Y(CO0_0_i));
    SLE bit_align_start (.D(N_1439_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        bit_align_done_0_sqmuxa_3_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        bit_align_start_Z));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_5 (.A(
        un10_tapcnt_final_5), .B(early_late_diff_Z[5]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_4_Z), .S(
        un1_early_late_diff_cry_5_S), .Y(un1_early_late_diff_cry_5_Y), 
        .FCO(un1_early_late_diff_cry_5_Z));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_66 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[6]), .C(un10_early_flags_2_Z[10]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[66]));
    SLE \late_flags[73]  (.D(late_flags_7_fast_Z[73]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[73]));
    SLE \early_flags[23]  (.D(early_flags_7_fast_Z[23]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[23]));
    CFG4 #( .INIT(16'h0B08) )  \tapcnt_final_13[4]  (.A(
        tapcnt_final_Z[4]), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .D(tapcnt_final_13_m1[4]), .Y(
        tapcnt_final_13_Z[4]));
    SLE \rst_cnt[0]  (.D(rst_cnt_s[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[0]));
    SLE \late_val[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[3])
        );
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_6 (.A(
        late_flags_pmux_126_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[57]), .D(late_flags_Z[121]), .FCI(
        late_flags_pmux_126_1_1_co0_2), .S(
        late_flags_pmux_126_1_1_wmux_6_S), .Y(
        late_flags_pmux_126_1_1_y7), .FCO(
        late_flags_pmux_126_1_1_co1_2));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_7 (.A(
        un16_tapcnt_final_7), .B(early_late_diff_Z[7]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_6_Z), .S(
        un1_early_late_diff_1_cry_7_S), .Y(
        un1_early_late_diff_1_cry_7_Y), .FCO(
        un1_early_late_diff_1_cry_7_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[17]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[17]), .C(
        un10_early_flags[17]), .Y(early_flags_7_fast_Z[17]));
    ARI1 #( .INIT(20'h472D8) )  \tap_cnt_RNO_0[6]  (.A(
        un1_tap_cnt_0_sqmuxa_14_0_Z[1]), .B(N_60), .C(tap_cnt_Z[6]), 
        .D(tapcnt_final_Z[6]), .FCI(tap_cnt_17_i_m2_cry_5), .S(N_74), 
        .Y(tap_cnt_RNO_0_Y[6]), .FCO(tap_cnt_RNO_0_FCO[6]));
    CFG3 #( .INIT(8'h04) )  early_last_set_2_sqmuxa (.A(
        restart_trng_fg_i), .B(early_val_0_sqmuxa_1_0_Z), .C(
        early_flags_pmux), .Y(early_last_set_2_sqmuxa_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_10 (.A(
        early_flags_pmux_63_1_0_0_y21), .B(
        early_flags_pmux_63_1_0_0_y9), .C(emflag_cnt_Z[2]), .D(VCC), 
        .FCI(early_flags_pmux_63_1_0_co0_4), .S(
        early_flags_pmux_63_1_0_wmux_10_S), .Y(
        early_flags_pmux_63_1_0_wmux_10_Y), .FCO(
        early_flags_pmux_63_1_0_co1_4));
    CFG4 #( .INIT(16'h0001) )  calc_done25_144 (.A(late_flags_Z[63]), 
        .B(late_flags_Z[62]), .C(late_flags_Z[61]), .D(
        late_flags_Z[60]), .Y(calc_done25_144_Z));
    CFG4 #( .INIT(16'h0007) )  rx_BIT_ALGN_MOVE_0_sqmuxa_2_1 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(
        rx_BIT_ALGN_MOVE_0_sqmuxa_0_Z), .C(
        un1_early_flags_1_sqmuxa_1_Z), .D(
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), .Y(
        rx_BIT_ALGN_MOVE_0_sqmuxa_2_1_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[119]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[119]), .C(
        un10_early_flags[119]), .Y(early_flags_7_fast_Z[119]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[4]  (.A(VCC), .B(
        rst_cnt_Z[4]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[3]), .S(
        rst_cnt_s[4]), .Y(rst_cnt_cry_Y_0[4]), .FCO(rst_cnt_cry_Z[4]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_19 (.A(
        early_flags_pmux_126_1_1_y7_0), .B(
        early_flags_pmux_126_1_1_y5_0), .C(emflag_cnt_Z[4]), .D(
        emflag_cnt_Z[3]), .FCI(early_flags_pmux_126_1_1_co1_8), .S(
        early_flags_pmux_126_1_1_wmux_19_S), .Y(
        early_flags_pmux_126_1_1_y0_8), .FCO(
        early_flags_pmux_126_1_1_co0_9));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_2 (.A(
        early_flags_pmux_126_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[51]), .D(early_flags_Z[115]), .FCI(
        early_flags_pmux_126_1_0_co0_0), .S(
        early_flags_pmux_126_1_0_wmux_2_S), .Y(
        early_flags_pmux_126_1_0_0_y3), .FCO(
        early_flags_pmux_126_1_0_co1_0));
    CFG4 #( .INIT(16'h8000) )  calc_done25_230 (.A(calc_done25_155_Z), 
        .B(calc_done25_154_Z), .C(calc_done25_153_Z), .D(
        calc_done25_152_Z), .Y(calc_done25_230_Z));
    SLE \late_flags[33]  (.D(late_flags_7_fast_Z[33]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[33]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[93]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[93]), .C(
        un10_early_flags[93]), .Y(early_flags_7_fast_Z[93]));
    SLE \early_flags[72]  (.D(early_flags_7_fast_Z[72]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[72]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[38]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[38]), .C(
        un10_early_flags[38]), .Y(late_flags_7_fast_Z[38]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_78 (.A(
        un10_early_flags_1_Z[72]), .B(un10_early_flags_1_Z[6]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_3_Z[46]), .Y(
        un10_early_flags[78]));
    SLE \bitalign_curr_state[1]  (.D(bitalign_curr_state_34[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[13]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[13]), .C(
        un10_early_flags[13]), .Y(late_flags_7_fast_Z[13]));
    SLE \late_flags[91]  (.D(late_flags_7_fast_Z[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[91]));
    SLE \restart_edge_reg[0]  (.D(Restart_trng_edge_det_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_edge_reg_Z[0]));
    SLE \early_flags[95]  (.D(early_flags_7_fast_Z[95]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[95]));
    CFG4 #( .INIT(16'h5150) )  rx_BIT_ALGN_LOAD_9_iv (.A(
        restart_trng_fg_i), .B(rx_err_Z), .C(un1_tap_cnt_0_sqmuxa_6_0), 
        .D(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z), .Y(rx_BIT_ALGN_LOAD_9)
        );
    SLE \rst_cnt[4]  (.D(rst_cnt_s[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[4]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[78]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[78]), .C(
        un10_early_flags[78]), .Y(early_flags_7_fast_Z[78]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[28]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[28]), .C(
        un10_early_flags[28]), .Y(late_flags_7_fast_Z[28]));
    CFG2 #( .INIT(4'h2) )  bitalign_curr_state154 (.A(
        bitalign_curr_state154_3_Z), .B(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state154_Z));
    CFG4 #( .INIT(16'h00CD) )  \bitalign_curr_state_34_4_0_.m67  (.A(
        m67_1), .B(m66_1), .C(bitalign_curr_state_Z[3]), .D(
        restart_trng_fg_i), .Y(bitalign_curr_state_34[1]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_184 (.A(early_flags_Z[23]), 
        .B(early_flags_Z[22]), .C(early_flags_Z[21]), .D(
        early_flags_Z[20]), .Y(calc_done25_184_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[123]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[123]), .C(
        un10_early_flags[123]), .Y(late_flags_7_fast_Z[123]));
    SLE \emflag_cnt[6]  (.D(emflag_cnt_s_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[6]));
    SLE \late_flags[120]  (.D(late_flags_7_fast_Z[120]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[120]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_76_2_0 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[5]), .Y(
        un10_early_flags_2_0[76]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[75]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[75]), .C(
        un10_early_flags[75]), .Y(early_flags_7_fast_Z[75]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_134 (.A(late_flags_Z[111]), 
        .B(late_flags_Z[110]), .C(late_flags_Z[109]), .D(
        late_flags_Z[108]), .Y(calc_done25_134_Z));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_2 (.A(
        tapcnt_final_upd_Z[2]), .B(tapcnt_final_Z[2]), .C(tap_cnt_Z[2])
        , .D(N_1416), .Y(bitalign_curr_state61_2_Z));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[6]  (.A(N_74), .B(N_63_0), .Y(
        N_1496_i));
    SLE \late_flags[8]  (.D(late_flags_7_fast_Z[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[8]));
    SLE \rst_cnt[2]  (.D(rst_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[2]));
    CFG3 #( .INIT(8'h20) )  rx_err_1_sqmuxa (.A(
        bitalign_curr_state162_Z), .B(un1_calc_done25_7_i), .C(
        early_flags_dec[127]), .Y(rx_err_1_sqmuxa_Z));
    SLE \no_early_no_late_val_end2[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[6]));
    SLE \early_flags[0]  (.D(early_flags_7_fast_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[0]));
    SLE calc_done (.D(N_1431_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(calc_done_0_sqmuxa_2_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(calc_done_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_158 (.A(late_flags_Z[15]), 
        .B(late_flags_Z[14]), .C(late_flags_Z[13]), .D(
        late_flags_Z[12]), .Y(calc_done25_158_Z));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_83 (.A(
        un10_early_flags_1_Z[80]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[0]), .Y(
        un10_early_flags[83]));
    SLE \early_flags[110]  (.D(early_flags_7_fast_Z[110]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[110]));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[5]  (.A(N_75), .B(N_63_0), .Y(
        N_1497_i));
    SLE \noearly_nolate_diff_nxt[2]  (.D(noearly_nolate_diff_nxt_8[2]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_2));
    CFG4 #( .INIT(16'h44F4) )  un1_bitalign_curr_state148_8_0 (.A(
        bit_align_dly_done_Z), .B(bitalign_curr_state163_Z), .C(
        bitalign_curr_state154_Z), .D(calc_done_0_sqmuxa_Z), .Y(
        un1_bitalign_curr_state148_8_0_Z));
    SLE \no_early_no_late_val_end1[2]  (.D(emflag_cnt_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[2]));
    SLE \no_early_no_late_val_end2[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[48]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[48]), .C(
        un10_early_flags[48]), .Y(late_flags_7_fast_Z[48]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_12 (.A(
        early_flags_pmux_126_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[39]), .D(early_flags_Z[103]), .FCI(
        early_flags_pmux_126_1_0_co0_5), .S(
        early_flags_pmux_126_1_0_wmux_12_S), .Y(
        early_flags_pmux_126_1_0_y1_0), .FCO(
        early_flags_pmux_126_1_0_co1_5));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIR4921[1]  (.A(
        no_early_no_late_val_st1_Z[1]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[1]), .Y(
        un1_no_early_no_late_val_st1_1_1[1]));
    SLE \late_flags[29]  (.D(late_flags_7_fast_Z[29]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[29]));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_34_4_0_.m34  (.A(
        early_flags_pmux), .B(early_cur_set_Z), .Y(N_35));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_123 (.A(
        un10_early_flags_1_Z[24]), .B(tap_cnt_Z[2]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[96]), .Y(
        un10_early_flags[123]));
    SLE \no_early_no_late_val_st1[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[81]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[81]), .C(
        un10_early_flags[81]), .Y(late_flags_7_fast_Z[81]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[119]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[119]), .C(
        un10_early_flags[119]), .Y(late_flags_7_fast_Z[119]));
    ARI1 #( .INIT(20'h4B4AA) )  \tapcnt_final_13_RNO[6]  (.A(
        un1_bitalign_curr_state169_12_sn), .B(early_val_Z[6]), .C(
        tapcnt_final_3_sqmuxa_Z), .D(tapcnt_final_13_m1_axb_6_1), .FCI(
        tapcnt_final_13_m1_cry_5), .S(tapcnt_final_13_m1[6]), .Y(
        tapcnt_final_13_RNO_Y[6]), .FCO(tapcnt_final_13_RNO_FCO[6]));
    CFG2 #( .INIT(4'h8) )  early_val_0_sqmuxa_1_0 (.A(
        bitalign_curr_state160_Z), .B(early_cur_set_Z), .Y(
        early_val_0_sqmuxa_1_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[67]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[67]), .C(
        un10_early_flags[67]), .Y(late_flags_7_fast_Z[67]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_71 (.A(tap_cnt_Z[6]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[71]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[19]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[19]), .C(
        un10_early_flags[19]), .Y(early_flags_7_fast_Z[19]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_6 (.A(late_val_Z[6])
        , .B(early_val_Z[6]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_5_Z), .S(tapcnt_final27_cry_6_S), .Y(
        tapcnt_final27_cry_6_Y), .FCO(tapcnt_final27));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_39 (.A(
        un10_early_flags_2_0[32]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[36]), .Y(un10_early_flags[39]));
    SLE \early_flags[4]  (.D(early_flags_7_fast_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[4]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_226 (.A(calc_done25_139_Z), 
        .B(calc_done25_138_Z), .C(calc_done25_137_Z), .D(
        calc_done25_136_Z), .Y(calc_done25_226_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[36]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[36]), .C(
        un10_early_flags[36]), .Y(early_flags_7_fast_Z[36]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_171 (.A(early_flags_Z[91]), 
        .B(early_flags_Z[90]), .C(early_flags_Z[89]), .D(
        early_flags_Z[88]), .Y(calc_done25_171_Z));
    SLE \late_flags[79]  (.D(late_flags_7_fast_Z[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[79]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_2 (.A(
        un10_tapcnt_final_2), .B(early_late_diff_Z[2]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_1_Z), .S(
        un1_early_late_diff_cry_2_S), .Y(un1_early_late_diff_cry_2_Y), 
        .FCO(un1_early_late_diff_cry_2_Z));
    CFG4 #( .INIT(16'hC0AC) )  un1_bitalign_curr_state148_2 (.A(
        bitalign_curr_state152_1_Z), .B(N_117_mux_1), .C(
        bitalign_curr_state_Z[3]), .D(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state148_2_Z));
    SLE \no_early_no_late_val_end2[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[1]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_1 (.A(
        un10_tapcnt_final_1), .B(early_late_diff_Z[1]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_0_Z), .S(
        un1_early_late_diff_cry_1_S), .Y(un1_early_late_diff_cry_1_Y), 
        .FCO(un1_early_late_diff_cry_1_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_0_0_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[2]), 
        .D(early_flags_Z[66]), .FCI(VCC), .S(
        early_flags_pmux_63_1_0_0_wmux_S), .Y(
        early_flags_pmux_63_1_0_0_y0), .FCO(
        early_flags_pmux_63_1_0_0_co0));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_0_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(un10_early_flags_2_0[0])
        );
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[40]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[40]), .C(
        un10_early_flags[40]), .Y(early_flags_7_fast_Z[40]));
    CFG4 #( .INIT(16'hFFFE) )  un1_bitalign_curr_state_1_sqmuxa_6 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_1_Z), .B(
        early_flags_0_sqmuxa_Z), .C(bitalign_curr_state_1_sqmuxa_4_Z), 
        .D(bit_align_done_0_sqmuxa_2_Z), .Y(
        un1_bitalign_curr_state_1_sqmuxa_6_i_0));
    CFG4 #( .INIT(16'hEA00) )  tapcnt_final_1_sqmuxa_2 (.A(
        calc_done26_Z), .B(calc_done27_Z), .C(
        un10_tapcnt_final_cry_7_Z), .D(bitalign_curr_state162_Z), .Y(
        tapcnt_final_1_sqmuxa_2_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_29 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_2_0[28]), .C(
        un10_early_flags_1_Z[5]), .Y(un10_early_flags[29]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[7]  (.A(VCC), .B(
        rst_cnt_Z[7]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[6]), .S(
        rst_cnt_s[7]), .Y(rst_cnt_cry_Y_0[7]), .FCO(rst_cnt_cry_Z[7]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[0]), .D(
        late_flags_Z[64]), .FCI(VCC), .S(late_flags_pmux_63_1_1_wmux_S)
        , .Y(late_flags_pmux_63_1_1_y0), .FCO(
        late_flags_pmux_63_1_1_co0));
    CFG3 #( .INIT(8'h80) )  bitalign_curr_state_0_sqmuxa_9 (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state155_Z), 
        .C(bitalign_curr_state61), .Y(bitalign_curr_state_0_sqmuxa_9_Z)
        );
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_1_wmux_8 (.A(
        early_flags_pmux_63_1_1_y0_3), .B(early_flags_pmux_63_1_1_y3), 
        .C(early_flags_pmux_63_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co0_3), .S(
        early_flags_pmux_63_1_1_wmux_8_S), .Y(
        early_flags_pmux_63_1_1_y9), .FCO(
        early_flags_pmux_63_1_1_co1_3));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_19 (.A(
        late_flags_pmux_63_1_1_y7_0), .B(late_flags_pmux_63_1_1_y5_0), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_63_1_1_co1_8), .S(
        late_flags_pmux_63_1_1_wmux_19_S), .Y(
        late_flags_pmux_63_1_1_y0_8), .FCO(
        late_flags_pmux_63_1_1_co0_9));
    CFG2 #( .INIT(4'h4) )  calc_done26 (.A(calc_done25_Z), .B(
        un1_tapcnt_final_Z), .Y(calc_done26_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[19]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[19]), .C(
        un10_early_flags[19]), .Y(late_flags_7_fast_Z[19]));
    SLE \late_flags[39]  (.D(late_flags_7_fast_Z[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[39]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_7 (.A(tap_cnt_Z[3]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[7]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_70 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_1_Z[64]), .C(
        un10_early_flags_2_0[64]), .Y(un10_early_flags[70]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIT6921[2]  (.A(
        no_early_no_late_val_st1_Z[2]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[2]), .Y(
        un1_no_early_no_late_val_st1_1_1[2]));
    SLE \late_flags[88]  (.D(late_flags_7_fast_Z[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[88]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_16_1 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[16]));
    SLE \late_flags[52]  (.D(late_flags_7_fast_Z[52]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[52]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_152 (.A(late_flags_Z[23]), 
        .B(late_flags_Z[22]), .C(late_flags_Z[21]), .D(
        late_flags_Z[20]), .Y(calc_done25_152_Z));
    CFG4 #( .INIT(16'hCC5F) )  \bitalign_curr_state_34_4_0_.m99  (.A(
        N_117_mux_1), .B(N_83), .C(rx_trng_done_Z), .D(
        bitalign_curr_state_Z[2]), .Y(N_100_0));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_6 (.A(
        un16_tapcnt_final_6), .B(early_late_diff_Z[6]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_5_Z), .S(
        un1_early_late_diff_1_cry_6_S), .Y(
        un1_early_late_diff_1_cry_6_Y), .FCO(
        un1_early_late_diff_1_cry_6_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[54]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[54]), .C(
        un10_early_flags[54]), .Y(early_flags_7_fast_Z[54]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_5_0 (.A(
        emflag_cnt_Z[5]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[5]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_4), .S(
        noearly_nolate_diff_nxt_8[5]), .Y(
        noearly_nolate_diff_nxt_8_cry_5_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_5));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_2 (.A(
        un10_tapcnt_final_2), .B(un16_tapcnt_final_2), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_1_Z), .S(
        un10_tapcnt_final_cry_2_S), .Y(un10_tapcnt_final_cry_2_Y), 
        .FCO(un10_tapcnt_final_cry_2_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_36_1 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[36]));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_2_0 (.A(
        emflag_cnt_Z[2]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[2]), .D(GND), .FCI(early_late_diff_8_cry_1), .S(
        early_late_diff_8[2]), .Y(early_late_diff_8_cry_2_0_Y), .FCO(
        early_late_diff_8_cry_2));
    SLE \late_flags[104]  (.D(late_flags_7_fast_Z[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[104]));
    SLE \early_flags[122]  (.D(early_flags_7_fast_Z[122]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[122]));
    SLE bit_align_dly_done (.D(bit_align_dly_done_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        bit_align_dly_done_0_sqmuxa_1_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bit_align_dly_done_Z));
    SLE \late_flags[0]  (.D(late_flags_7_fast_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[0]));
    SLE \restart_reg[1]  (.D(restart_reg_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_reg_Z[1]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_6_0 (
        .A(emflag_cnt_Z[6]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[6]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_5), .S(
        noearly_nolate_diff_start_7[6]), .Y(
        noearly_nolate_diff_start_7_cry_6_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_6));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_13 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[3]), .C(un10_early_flags_1_Z[5]), .D(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[13]));
    SLE \late_flags[18]  (.D(late_flags_7_fast_Z[18]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[18]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_4 (.A(
        late_flags_pmux_63_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[40]), .D(late_flags_Z[104]), .FCI(
        late_flags_pmux_63_1_1_co0_1), .S(
        late_flags_pmux_63_1_1_wmux_4_S), .Y(late_flags_pmux_63_1_1_y5)
        , .FCO(late_flags_pmux_63_1_1_co1_1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[83]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[83]), .C(
        un10_early_flags[83]), .Y(late_flags_7_fast_Z[83]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[116]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[116]), .C(
        un10_early_flags[116]), .Y(early_flags_7_fast_Z[116]));
    CFG2 #( .INIT(4'h1) )  bitalign_curr_state148_2 (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[4]), .Y(
        bitalign_curr_state148_2_Z));
    CFG4 #( .INIT(16'hCCDF) )  rx_err_0_sqmuxa_1_i (.A(
        bitalign_curr_state162_Z), .B(restart_trng_fg_i), .C(
        un1_calc_done25_7_i), .D(un1_bitalign_curr_state148_9_2_Z), .Y(
        rx_err_0_sqmuxa_1_i_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[73]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[73]), .C(
        un10_early_flags[73]), .Y(early_flags_7_fast_Z[73]));
    CFG2 #( .INIT(4'hE) )  \un1_tap_cnt_0_sqmuxa_14_0_o2_0[1]  (.A(
        un1_bitalign_curr_state_1_sqmuxa_2_i_0), .B(
        rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), .Y(N_82));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_1_0 (
        .A(emflag_cnt_Z[1]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[1]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_0), .S(
        noearly_nolate_diff_start_7[1]), .Y(
        noearly_nolate_diff_start_7_cry_1_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_1));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_6 (.A(
        early_flags_pmux_63_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[58]), .D(early_flags_Z[122]), .FCI(
        early_flags_pmux_63_1_0_co0_2), .S(
        early_flags_pmux_63_1_0_wmux_6_S), .Y(
        early_flags_pmux_63_1_0_0_y7), .FCO(
        early_flags_pmux_63_1_0_co1_2));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_0_wmux_9 (.A(VCC), 
        .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_63_1_0_co1_3), .S(
        late_flags_pmux_63_1_0_wmux_9_S), .Y(
        late_flags_pmux_63_1_0_wmux_9_Y), .FCO(
        late_flags_pmux_63_1_0_co0_4));
    SLE \early_flags[54]  (.D(early_flags_7_fast_Z[54]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[54]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_4 (.A(
        un16_tapcnt_final_4), .B(un10_tapcnt_final_4), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_3_Z), .S(
        un16_tapcnt_final_cry_4_S), .Y(un16_tapcnt_final_cry_4_Y), 
        .FCO(un16_tapcnt_final_cry_4_Z));
    CFG4 #( .INIT(16'hFFFD) )  un1_bitalign_curr_state148_9_2 (.A(
        un1_bitalign_curr_state148_5_Z), .B(
        un1_bitalign_curr_state148_9_0_Z), .C(early_flags_1_sqmuxa_1_Z)
        , .D(early_flags_0_sqmuxa_1_Z), .Y(
        un1_bitalign_curr_state148_9_2_Z));
    SLE \early_flags[43]  (.D(early_flags_7_fast_Z[43]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[43]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[44]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[44]), .C(
        un10_early_flags[44]), .Y(early_flags_7_fast_Z[44]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_233 (.A(calc_done25_167_Z), 
        .B(calc_done25_166_Z), .C(calc_done25_165_Z), .D(
        calc_done25_164_Z), .Y(calc_done25_233_Z));
    SLE \late_flags[48]  (.D(late_flags_7_fast_Z[48]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[48]));
    SLE \late_flags[62]  (.D(late_flags_7_fast_Z[62]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[62]));
    CFG4 #( .INIT(16'h083B) )  \bitalign_curr_state_34_4_0_.m86_1  (.A(
        bitalign_curr_state161_2_Z), .B(bitalign_curr_state_Z[4]), .C(
        N_76_0), .D(N_75_0), .Y(m86_1));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[16]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[16]), .C(
        un10_early_flags[16]), .Y(late_flags_7_fast_Z[16]));
    SLE \late_flags[123]  (.D(late_flags_7_fast_Z[123]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[123]));
    SLE \late_flags[109]  (.D(late_flags_7_fast_Z[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[109]));
    SLE \early_late_diff[3]  (.D(early_late_diff_8[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[3]));
    CFG4 #( .INIT(16'h4C7F) )  \bitalign_curr_state_34_4_0_.m101_1_1  
        (.A(bitalign_curr_state161_2_Z), .B(bitalign_curr_state_Z[4]), 
        .C(N_94), .D(N_92), .Y(m101_1_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[109]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[109]), .C(
        un10_early_flags[109]), .Y(early_flags_7_fast_Z[109]));
    SLE \early_late_diff[6]  (.D(early_late_diff_8[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[6]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_156 (.A(late_flags_Z[7]), 
        .B(late_flags_Z[6]), .C(late_flags_Z[5]), .D(late_flags_Z[4]), 
        .Y(calc_done25_156_Z));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_1 (.A(
        tapcnt_final_upd_Z[1]), .B(tapcnt_final_Z[1]), .C(tap_cnt_Z[1])
        , .D(N_1416), .Y(bitalign_curr_state61_1_Z));
    CFG2 #( .INIT(4'h4) )  \bitalign_curr_state_RNISUK8[0]  (.A(
        bitalign_curr_state_Z[0]), .B(bitalign_curr_state_Z[2]), .Y(
        N_1456_1));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_0_wmux_16 (.A(
        early_flags_pmux_126_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[47]), .D(early_flags_Z[111]), .FCI(
        early_flags_pmux_126_1_0_co0_7), .S(
        early_flags_pmux_126_1_0_wmux_16_S), .Y(
        early_flags_pmux_126_1_0_y5_0), .FCO(
        early_flags_pmux_126_1_0_co1_7));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_111 (.A(
        un10_early_flags_1_Z[96]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[111]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[91]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[91]), .C(
        un10_early_flags[91]), .Y(late_flags_7_fast_Z[91]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNI0M2N6[1]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIJGIR_Z[1]), .B(
        early_val_RNI6O2D1_Z[1]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[1]), .FCI(tapcnt_final_13_m1_cry_0), .S(
        tapcnt_final_13_m1[1]), .Y(early_val_RNI0M2N6_Y[1]), .FCO(
        tapcnt_final_13_m1_cry_1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[115]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[115]), .C(
        un10_early_flags[115]), .Y(early_flags_7_fast_Z[115]));
    CFG4 #( .INIT(16'h10BA) )  \bitalign_curr_state_34_4_0_.m82_1_1  (
        .A(bitalign_curr_state_Z[1]), .B(early_flags_dec[127]), .C(
        bitalign_curr_state89_Z), .D(N_63), .Y(m82_1_1));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_6 (.A(
        late_flags_pmux_63_1_0_y0_2), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[58]), .D(late_flags_Z[122]), .FCI(
        late_flags_pmux_63_1_0_co0_2), .S(
        late_flags_pmux_63_1_0_wmux_6_S), .Y(
        late_flags_pmux_63_1_0_0_y7), .FCO(
        late_flags_pmux_63_1_0_co1_2));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNII43D1[5]  (.A(early_val_Z[5])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[5]), .Y(
        early_val_RNII43D1_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[100]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[100]), .C(
        un10_early_flags[100]), .Y(late_flags_7_fast_Z[100]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[114]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[114]), .C(
        un10_early_flags[114]), .Y(early_flags_7_fast_Z[114]));
    CFG3 #( .INIT(8'h01) )  bit_align_done_0_sqmuxa_3_1 (.A(
        bitalign_curr_state_1_sqmuxa_4_Z), .B(restart_trng_fg_i), .C(
        bit_align_dly_done_0_sqmuxa_Z), .Y(
        bit_align_done_0_sqmuxa_3_1_Z));
    CFG4 #( .INIT(16'h0002) )  un1_tapcnt_final_0_sqmuxa_RNO (.A(
        calc_done_4_sqmuxa_0_Z), .B(un1_calc_done25_5_Z), .C(
        tapcnt_final27), .D(restart_trng_fg_i), .Y(
        tapcnt_final_5_sqmuxa));
    SLE \late_flags[121]  (.D(late_flags_7_fast_Z[121]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[121]));
    CFG4 #( .INIT(16'h0004) )  calc_done28 (.A(un1_tapcnt_final_Z), .B(
        un1_noearly_nolate_diff_nxt_valid_Z), .C(calc_done25_Z), .D(
        un1_noearly_nolate_diff_start_valid_Z), .Y(calc_done28_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[5]  (.A(VCC), .B(
        rst_cnt_Z[5]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[4]), .S(
        rst_cnt_s[5]), .Y(rst_cnt_cry_Y_0[5]), .FCO(rst_cnt_cry_Z[5]));
    SLE \tapcnt_final_upd[2]  (.D(tapcnt_final_upd_8_cry_2_0_Y), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[2]));
    SLE sig_rx_BIT_ALGN_CLR_FLGS (.D(sig_rx_BIT_ALGN_CLR_FLGS_11), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_2_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(sig_rx_BIT_ALGN_CLR_FLGS_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_63_1_0_co1_3), .S(
        early_flags_pmux_63_1_0_wmux_9_S), .Y(
        early_flags_pmux_63_1_0_wmux_9_Y), .FCO(
        early_flags_pmux_63_1_0_co0_4));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_10 (.A(
        early_flags_pmux_126_1_1_y21), .B(early_flags_pmux_126_1_1_y9), 
        .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_126_1_1_co0_4), .S(
        early_flags_pmux_126_1_1_wmux_10_S), .Y(
        early_flags_pmux_126_1_1_wmux_10_Y), .FCO(
        early_flags_pmux_126_1_1_co1_4));
    CFG4 #( .INIT(16'h3A00) )  \bitalign_curr_state_34_4_0_.m106  (.A(
        N_108), .B(N_63), .C(bitalign_curr_state_Z[1]), .D(i22_mux_1), 
        .Y(i22_mux));
    CFG4 #( .INIT(16'hFFFE) )  emflag_cnt_1_sqmuxa_1_RNIGA491 (.A(
        emflag_cnt_1_sqmuxa_1_Z), .B(bitalign_curr_state_1_sqmuxa_4_Z), 
        .C(tap_cnt_0_sqmuxa_1_Z), .D(emflag_cntlde_1), .Y(
        emflag_cntlde_4));
    CFG3 #( .INIT(8'hFE) )  un1_tapcnt_final_0_sqmuxa (.A(
        tapcnt_final_5_sqmuxa), .B(un1_bitalign_curr_state_12_Z), .C(
        un1_restart_trng_fg_10_sn), .Y(un1_tapcnt_final_0_sqmuxa_Z));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_s[9]  (.A(VCC), .B(
        rst_cnt_Z[9]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[8]), .S(
        rst_cnt_s_Z[9]), .Y(rst_cnt_s_Y_0[9]), .FCO(rst_cnt_s_FCO_0[9])
        );
    SLE \late_flags[84]  (.D(late_flags_7_fast_Z[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[84]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[117]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[117]), .C(
        un10_early_flags[117]), .Y(late_flags_7_fast_Z[117]));
    SLE \late_val[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[4])
        );
    SLE \early_flags[56]  (.D(early_flags_7_fast_Z[56]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[56]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[60]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[60]), .C(
        un10_early_flags[60]), .Y(late_flags_7_fast_Z[60]));
    SLE \early_flags[57]  (.D(early_flags_7_fast_Z[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[57]));
    CFG3 #( .INIT(8'h20) )  bitalign_curr_state149 (.A(N_117_mux_1), 
        .B(bitalign_curr_state_Z[4]), .C(i22_mux_1), .Y(
        bitalign_curr_state149_Z));
    CFG4 #( .INIT(16'h00A8) )  calc_done_RNO (.A(
        bitalign_curr_state_Z[4]), .B(early_flags_dec[127]), .C(
        un1_calc_done25_7_i), .D(restart_trng_fg_i), .Y(N_1431_i));
    CFG3 #( .INIT(8'h8B) )  \early_val_RNI9R2D1[2]  (.A(early_val_Z[2])
        , .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_st1_1_1[2]), .Y(
        early_val_RNI9R2D1_Z[2]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_18 (.A(
        early_flags_pmux_63_1_1_y0_7), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[60]), .D(early_flags_Z[124]), .FCI(
        early_flags_pmux_63_1_1_co0_8), .S(
        early_flags_pmux_63_1_1_wmux_18_S), .Y(
        early_flags_pmux_63_1_1_y7_0), .FCO(
        early_flags_pmux_63_1_1_co1_8));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_12 (.A(
        late_flags_pmux_126_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[39]), .D(late_flags_Z[103]), .FCI(
        late_flags_pmux_126_1_0_co0_5), .S(
        late_flags_pmux_126_1_0_wmux_12_S), .Y(
        late_flags_pmux_126_1_0_y1_0), .FCO(
        late_flags_pmux_126_1_0_co1_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[105]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[105]), .C(
        un10_early_flags[105]), .Y(late_flags_7_fast_Z[105]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[13]), 
        .D(early_flags_Z[77]), .FCI(early_flags_pmux_126_1_1_co1_6), 
        .S(early_flags_pmux_126_1_1_wmux_15_S), .Y(
        early_flags_pmux_126_1_1_y0_6), .FCO(
        early_flags_pmux_126_1_1_co0_7));
    CFG4 #( .INIT(16'h4000) )  bitalign_curr_state163 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state163_2), .D(bitalign_curr_state_Z[1]), .Y(
        bitalign_curr_state163_Z));
    CFG3 #( .INIT(8'hFE) )  early_flags_1_sqmuxa_RNIRGCS (.A(
        early_flags_1_sqmuxa_Z), .B(un1_tap_cnt_0_sqmuxa_6_0), .C(
        restart_trng_fg_i), .Y(early_flags_0_sqmuxa_2_i));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_2 (.A(
        late_flags_pmux_126_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[51]), .D(late_flags_Z[115]), .FCI(
        late_flags_pmux_126_1_0_co0_0), .S(
        late_flags_pmux_126_1_0_wmux_2_S), .Y(
        late_flags_pmux_126_1_0_0_y3), .FCO(
        late_flags_pmux_126_1_0_co1_0));
    CFG2 #( .INIT(4'h8) )  early_flags_0_sqmuxa (.A(
        bitalign_curr_state153_Z), .B(BIT_ALGN_OOR_c), .Y(
        early_flags_0_sqmuxa_Z));
    SLE \late_flags[14]  (.D(late_flags_7_fast_Z[14]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[14]));
    SLE \early_flags[51]  (.D(early_flags_7_fast_Z[51]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[51]));
    SLE \early_flags[10]  (.D(early_flags_7_fast_Z[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[10]));
    ARI1 #( .INIT(20'h572D8) )  \tapcnt_final_RNIOTM22[1]  (.A(
        un1_tap_cnt_0_sqmuxa_14_0_Z[1]), .B(N_60), .C(tap_cnt_Z[1]), 
        .D(tapcnt_final_Z[1]), .FCI(tap_cnt_17_i_m2_cry_0), .S(N_79), 
        .Y(tapcnt_final_RNIOTM22_Y[1]), .FCO(tap_cnt_17_i_m2_cry_1));
    SLE \no_early_no_late_val_st2[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[0]));
    SLE mv_dn_fg (.D(tapcnt_final_upd_3_sqmuxa_1), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(mv_dn_fg_0_sqmuxa_i_0_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(mv_dn_fg_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_72_1 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_1_Z[72]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_178 (.A(early_flags_Z[63]), 
        .B(early_flags_Z[62]), .C(early_flags_Z[61]), .D(
        early_flags_Z[60]), .Y(calc_done25_178_Z));
    GND GND_Z (.Y(GND));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[11]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[11]), .C(
        un10_early_flags[11]), .Y(early_flags_7_fast_Z[11]));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_1 (.A(
        un16_tapcnt_final_1), .B(un10_tapcnt_final_1), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_0_Z), .S(
        un16_tapcnt_final_cry_1_S), .Y(un16_tapcnt_final_cry_1_Y), 
        .FCO(un16_tapcnt_final_cry_1_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_16 (.A(
        late_flags_pmux_126_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[47]), .D(late_flags_Z[111]), .FCI(
        late_flags_pmux_126_1_0_co0_7), .S(
        late_flags_pmux_126_1_0_wmux_16_S), .Y(
        late_flags_pmux_126_1_0_y5_0), .FCO(
        late_flags_pmux_126_1_0_co1_7));
    SLE \early_flags[39]  (.D(early_flags_7_fast_Z[39]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[39]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_101 (.A(
        un10_early_flags_1_Z[96]), .B(un10_early_flags_1_Z[5]), .C(
        un10_early_flags_2_0[100]), .Y(un10_early_flags[101]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_191 (.A(early_flags_Z[11]), 
        .B(early_flags_Z[10]), .C(early_flags_Z[9]), .D(
        early_flags_Z[8]), .Y(calc_done25_191_Z));
    SLE \no_early_no_late_val_st1[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[4]));
    SLE \late_flags[98]  (.D(late_flags_7_fast_Z[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[98]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_129 (.A(late_flags_Z[115]), 
        .B(late_flags_Z[114]), .C(late_flags_Z[113]), .D(
        late_flags_Z[112]), .Y(calc_done25_129_Z));
    SLE \late_val[5]  (.D(emflag_cnt_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[5])
        );
    SLE \late_flags[44]  (.D(late_flags_7_fast_Z[44]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[44]));
    CFG2 #( .INIT(4'h8) )  un1_retrain_adj_tap (.A(mv_up_fg_Z), .B(
        mv_dn_fg_Z), .Y(un1_retrain_adj_tap_i));
    CFG1 #( .INIT(2'h1) )  \rst_cnt_RNO[0]  (.A(rst_cnt_Z[0]), .Y(
        rst_cnt_s[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[55]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[55]), .C(
        un10_early_flags[55]), .Y(late_flags_7_fast_Z[55]));
    SLE \late_flags[105]  (.D(late_flags_7_fast_Z[105]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[105]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_16 (.A(
        late_flags_pmux_63_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[46]), .D(late_flags_Z[110]), .FCI(
        late_flags_pmux_63_1_0_co0_7), .S(
        late_flags_pmux_63_1_0_wmux_16_S), .Y(
        late_flags_pmux_63_1_0_y5_0), .FCO(
        late_flags_pmux_63_1_0_co1_7));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_125 (.A(tap_cnt_Z[1]), 
        .B(un10_early_flags_1_Z[5]), .C(un10_early_flags_1_Z[24]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[125]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_244 (.A(calc_done25_160_Z), 
        .B(calc_done25_161_Z), .C(calc_done25_233_Z), .D(
        calc_done25_209_Z), .Y(calc_done25_244_Z));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_126_1_1_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        late_flags_pmux_126_1_1_co1_3), .S(
        late_flags_pmux_126_1_1_wmux_9_S), .Y(
        late_flags_pmux_126_1_1_wmux_9_Y), .FCO(
        late_flags_pmux_126_1_1_co0_4));
    SLE \early_flags[8]  (.D(early_flags_7_fast_Z[8]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[8]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[89]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[89]), .C(
        un10_early_flags[89]), .Y(late_flags_7_fast_Z[89]));
    SLE \late_flags[112]  (.D(late_flags_7_fast_Z[112]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[112]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_40_2_0 (.A(tap_cnt_Z[2]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[40]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_44_2_0 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[4]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[44]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_12 (.A(
        early_flags_pmux_63_1_0_y0_4), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[38]), .D(early_flags_Z[102]), .FCI(
        early_flags_pmux_63_1_0_co0_5), .S(
        early_flags_pmux_63_1_0_wmux_12_S), .Y(
        early_flags_pmux_63_1_0_y1_0), .FCO(
        early_flags_pmux_63_1_0_co1_5));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_24_1 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[3]), .Y(un10_early_flags_1_Z[24]));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_4 (.A(
        early_flags_pmux_63_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[40]), .D(early_flags_Z[104]), .FCI(
        early_flags_pmux_63_1_1_co0_1), .S(
        early_flags_pmux_63_1_1_wmux_4_S), .Y(
        early_flags_pmux_63_1_1_y5), .FCO(
        early_flags_pmux_63_1_1_co1_1));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_15 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[15]), 
        .D(early_flags_Z[79]), .FCI(early_flags_pmux_126_1_0_co1_6), 
        .S(early_flags_pmux_126_1_0_wmux_15_S), .Y(
        early_flags_pmux_126_1_0_y0_6), .FCO(
        early_flags_pmux_126_1_0_co0_7));
    SLE \early_flags[84]  (.D(early_flags_7_fast_Z[84]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[84]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[4]), 
        .D(early_flags_Z[68]), .FCI(early_flags_pmux_63_1_1_co1_4), .S(
        early_flags_pmux_63_1_1_wmux_11_S), .Y(
        early_flags_pmux_63_1_1_y0_4), .FCO(
        early_flags_pmux_63_1_1_co0_5));
    CFG4 #( .INIT(16'hFE00) )  bitalign_curr_state12_0_0 (.A(
        BIT_ALGN_EYE_IN_c[2]), .B(BIT_ALGN_EYE_IN_c[1]), .C(
        BIT_ALGN_EYE_IN_c[0]), .D(PLL_LOCK_0), .Y(
        bitalign_curr_state12_0));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[26]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[26]), .C(
        un10_early_flags[26]), .Y(early_flags_7_fast_Z[26]));
    CFG3 #( .INIT(8'h01) )  un10_early_flags_28_2_0 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[1]), .C(tap_cnt_Z[6]), .Y(
        un10_early_flags_2_0[28]));
    CFG4 #( .INIT(16'hBBBA) )  \un1_tap_cnt_0_sqmuxa_14_0[1]  (.A(
        restart_trng_fg_i), .B(un1_early_flags_1_sqmuxa_i), .C(N_82), 
        .D(bitalign_curr_state_0_sqmuxa_10), .Y(
        un1_tap_cnt_0_sqmuxa_14_0_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[86]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[86]), .C(
        un10_early_flags[86]), .Y(early_flags_7_fast_Z[86]));
    SLE \early_flags[69]  (.D(early_flags_7_fast_Z[69]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[69]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[93]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[93]), .C(
        un10_early_flags[93]), .Y(late_flags_7_fast_Z[93]));
    SLE \early_flags[12]  (.D(early_flags_7_fast_Z[12]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[12]));
    CFG4 #( .INIT(16'hDFFF) )  \late_flags_7_i_o4[49]  (.A(
        tap_cnt_Z[0]), .B(tap_cnt_Z[1]), .C(un10_early_flags_2_0[48]), 
        .D(un10_early_flags_1_Z[48]), .Y(N_208));
    SLE \no_early_no_late_val_st2[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[3]));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_101_2 (.A(tap_cnt_Z[5]), 
        .B(tap_cnt_Z[6]), .Y(un10_early_flags_1_Z[96]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[26]), 
        .D(late_flags_Z[90]), .FCI(late_flags_pmux_63_1_0_co1_1), .S(
        late_flags_pmux_63_1_0_wmux_5_S), .Y(
        late_flags_pmux_63_1_0_y0_2), .FCO(
        late_flags_pmux_63_1_0_co0_2));
    CFG4 #( .INIT(16'h8000) )  calc_done25_234 (.A(calc_done25_171_Z), 
        .B(calc_done25_170_Z), .C(calc_done25_169_Z), .D(
        calc_done25_168_Z), .Y(calc_done25_234_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_48_1 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[4]), .Y(un10_early_flags_1_Z[48]));
    CFG2 #( .INIT(4'h7) )  un10_early_flags_18_1_i (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[1]), .Y(N_1499));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[120]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[120]), .C(
        un10_early_flags[120]), .Y(late_flags_7_fast_Z[120]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_0_wmux_7 (.A(
        early_flags_pmux_63_1_0_0_y7), .B(early_flags_pmux_63_1_0_0_y5)
        , .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_0_co1_2), .S(
        early_flags_pmux_63_1_0_wmux_7_S), .Y(
        early_flags_pmux_63_1_0_y0_3), .FCO(
        early_flags_pmux_63_1_0_co0_3));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_92 (.A(
        un10_early_flags_1_Z[12]), .B(un10_early_flags_1_Z[0]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_1_Z[80]), .Y(
        un10_early_flags[92]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[66]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[66]), .C(
        un10_early_flags[66]), .Y(early_flags_7_fast_Z[66]));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_start_7_s_7 (.A(
        VCC), .B(un1_restart_trng_fg_5_Z), .C(GND), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_6), .S(
        noearly_nolate_diff_start_7[7]), .Y(
        noearly_nolate_diff_start_7_s_7_Y), .FCO(
        noearly_nolate_diff_start_7_s_7_FCO));
    CFG2 #( .INIT(4'h8) )  tap_cnt_0_sqmuxa_1 (.A(
        bitalign_curr_state148_Z), .B(bitalign_curr_state12_Z), .Y(
        tap_cnt_0_sqmuxa_1_Z));
    SLE mv_up_fg (.D(tapcnt_final_upd_2_sqmuxa_1), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(mv_up_fg_0_sqmuxa_i_0_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(mv_up_fg_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_74 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_1_Z[10]), .C(
        un10_early_flags_2_0[72]), .Y(un10_early_flags[74]));
    SLE \late_flags[2]  (.D(late_flags_7_fast_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[2]));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI9ABM[0]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[0]), .D(GND), .FCI(
        timeout_cnt_cry_cy), .S(timeout_cnt_s[0]), .Y(
        timeout_cnt_RNI9ABM_Y[0]), .FCO(timeout_cnt_cry[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_4 (.A(
        late_flags_pmux_126_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[41]), .D(late_flags_Z[105]), .FCI(
        late_flags_pmux_126_1_1_co0_1), .S(
        late_flags_pmux_126_1_1_wmux_4_S), .Y(
        late_flags_pmux_126_1_1_y5), .FCO(
        late_flags_pmux_126_1_1_co1_1));
    SLE \early_flags[86]  (.D(early_flags_7_fast_Z[86]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[86]));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_start_7_cry_0_0_cy 
        (.A(VCC), .B(un1_restart_trng_fg_5_Z), .C(GND), .D(GND), .FCI(
        VCC), .S(noearly_nolate_diff_start_7_cry_0_0_cy_S), .Y(
        noearly_nolate_diff_start_7_cry_0_0_cy_Y), .FCO(
        noearly_nolate_diff_start_7_cry_0_0_cy_Z));
    SLE \early_flags[9]  (.D(early_flags_7_fast_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[9]));
    SLE \early_flags[94]  (.D(early_flags_7_fast_Z[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[94]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_172 (.A(early_flags_Z[71]), 
        .B(early_flags_Z[70]), .C(early_flags_Z[69]), .D(
        early_flags_Z[68]), .Y(calc_done25_172_Z));
    CFG4 #( .INIT(16'h1000) )  un10_early_flags_113 (.A(tap_cnt_Z[3]), 
        .B(N_1498), .C(un10_early_flags_2_Z[8]), .D(
        un10_early_flags_1_Z[96]), .Y(un10_early_flags[113]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[75]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[75]), .C(
        un10_early_flags[75]), .Y(late_flags_7_fast_Z[75]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[86]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[86]), .C(
        un10_early_flags[86]), .Y(late_flags_7_fast_Z[86]));
    SLE \early_flags[87]  (.D(early_flags_7_fast_Z[87]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[87]));
    SLE \late_flags[127]  (.D(late_flags_7_fast_Z[127]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[127]));
    ARI1 #( .INIT(20'h0EC2C) )  late_flags_pmux_63_1_1_wmux_10 (.A(
        late_flags_pmux_63_1_1_y21), .B(late_flags_pmux_63_1_1_y9), .C(
        emflag_cnt_Z[2]), .D(VCC), .FCI(late_flags_pmux_63_1_1_co0_4), 
        .S(late_flags_pmux_63_1_1_wmux_10_S), .Y(
        late_flags_pmux_63_1_1_wmux_10_Y), .FCO(
        late_flags_pmux_63_1_1_co1_4));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[125]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[125]), .C(
        un10_early_flags[125]), .Y(late_flags_7_fast_Z[125]));
    SLE rx_trng_done (.D(N_1403), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(rx_trng_done_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(rx_trng_done_Z));
    SLE \late_flags[94]  (.D(late_flags_7_fast_Z[94]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[94]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[68]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[68]), .C(
        un10_early_flags[68]), .Y(late_flags_7_fast_Z[68]));
    SLE \early_flags[81]  (.D(early_flags_7_fast_Z[81]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[81]));
    SLE late_cur_set (.D(late_cur_set_2_sqmuxa_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        late_cur_set_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(late_cur_set_Z));
    SLE \early_flags[79]  (.D(early_flags_7_fast_Z[79]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[79]));
    CFG4 #( .INIT(16'hFFFE) )  bitalign_curr_state61_NE_4 (.A(
        bitalign_curr_state61_6_Z), .B(bitalign_curr_state61_3_Z), .C(
        bitalign_curr_state61_2_Z), .D(bitalign_curr_state61_1_Z), .Y(
        bitalign_curr_state61_NE_4_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[106]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[106]), .C(
        un10_early_flags[106]), .Y(early_flags_7_fast_Z[106]));
    SLE \retrain_reg[2]  (.D(retrain_reg_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(retrain_reg_Z[2]));
    CFG2 #( .INIT(4'hD) )  \bitalign_curr_state_34_4_0_.m68  (.A(
        bitalign_curr_state13), .B(bitalign_curr_state_Z[0]), .Y(N_69));
    SLE \late_val[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[1])
        );
    CFG2 #( .INIT(4'h1) )  un10_early_flags_0_1 (.A(tap_cnt_Z[0]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_1_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[112]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[112]), .C(
        un10_early_flags[112]), .Y(early_flags_7_fast_Z[112]));
    SLE \early_flags[104]  (.D(early_flags_7_fast_Z[104]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[104]));
    SLE \emflag_cnt[3]  (.D(emflag_cnt_s[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[58]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[58]), .C(
        un10_early_flags[58]), .Y(early_flags_7_fast_Z[58]));
    ARI1 #( .INIT(20'h55104) )  tapcnt_final_upd_8_cry_2_0 (.A(
        tap_cnt_Z[2]), .B(mv_dn_fg_0_sqmuxa_i_o2_Z), .C(N_100), .D(
        mv_up_fg_Z), .FCI(GND), .S(tapcnt_final_upd_8_cry_2_0_S), .Y(
        tapcnt_final_upd_8_cry_2_0_Y), .FCO(tapcnt_final_upd_8_cry_2));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[1]  (.A(VCC), .B(
        rst_cnt_Z[1]), .C(GND), .D(GND), .FCI(rst_cnt_s_715_FCO), .S(
        rst_cnt_s[1]), .Y(rst_cnt_cry_Y_0[1]), .FCO(rst_cnt_cry_Z[1]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_21_2 (.A(tap_cnt_Z[4]), .B(
        tap_cnt_Z[1]), .Y(un10_early_flags_2_Z[21]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_154 (.A(late_flags_Z[31]), 
        .B(late_flags_Z[30]), .C(late_flags_Z[29]), .D(
        late_flags_Z[28]), .Y(calc_done25_154_Z));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_80_1 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[4]), .Y(un10_early_flags_1_Z[80]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_163 (.A(early_flags_Z[123]), 
        .B(early_flags_Z[122]), .C(early_flags_Z[121]), .D(
        early_flags_Z[120]), .Y(calc_done25_163_Z));
    SLE \no_early_no_late_val_end1[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[57]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[57]), .C(
        un10_early_flags[57]), .Y(late_flags_7_fast_Z[57]));
    ARI1 #( .INIT(20'h45500) )  early_late_diff_8_s_7 (.A(VCC), .B(
        un1_restart_trng_fg_5_Z), .C(GND), .D(GND), .FCI(
        early_late_diff_8_cry_6), .S(early_late_diff_8[7]), .Y(
        early_late_diff_8_s_7_Y), .FCO(early_late_diff_8_s_7_FCO));
    SLE \tapcnt_final_upd[5]  (.D(tapcnt_final_upd_8[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[5]));
    SLE \noearly_nolate_diff_start[5]  (.D(
        noearly_nolate_diff_start_7[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_5));
    SLE \early_flags[58]  (.D(early_flags_7_fast_Z[58]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[58]));
    CFG4 #( .INIT(16'h1300) )  \bitalign_curr_state_34_4_0_.m19  (.A(
        late_cur_set_Z), .B(early_cur_set_Z), .C(late_flags_pmux), .D(
        early_flags_pmux), .Y(N_20));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[55]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[55]), .C(
        un10_early_flags[55]), .Y(early_flags_7_fast_Z[55]));
    SLE \early_flags[96]  (.D(early_flags_7_fast_Z[96]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[96]));
    SLE \emflag_cnt[2]  (.D(emflag_cnt_s[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(emflag_cnte), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(emflag_cnt_Z[2]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[5]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[5]), .C(
        un10_early_flags[5]), .Y(early_flags_7_fast_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[16]), 
        .D(late_flags_Z[80]), .FCI(late_flags_pmux_63_1_1_co1), .S(
        late_flags_pmux_63_1_1_wmux_1_S), .Y(
        late_flags_pmux_63_1_1_y0_0), .FCO(
        late_flags_pmux_63_1_1_co0_0));
    SLE \early_flags[97]  (.D(early_flags_7_fast_Z[97]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[97]));
    SLE \early_flags[126]  (.D(early_flags_7_fast_Z[126]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[126]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_176 (.A(early_flags_Z[55]), 
        .B(early_flags_Z[54]), .C(early_flags_Z[53]), .D(
        early_flags_Z[52]), .Y(calc_done25_176_Z));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_4 (.A(
        tapcnt_final_upd_Z[4]), .B(tapcnt_final_Z[4]), .C(tap_cnt_Z[4])
        , .D(N_1416), .Y(bitalign_curr_state61_4_Z));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_64_1 (.A(tap_cnt_Z[6]), .B(
        tap_cnt_Z[0]), .Y(un10_early_flags_1_Z[64]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[101]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[101]), .C(
        un10_early_flags[101]), .Y(late_flags_7_fast_Z[101]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_103 (.A(
        un10_early_flags_1_Z[36]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[4]), .D(un10_early_flags_3_Z[87]), .Y(
        un10_early_flags[103]));
    CFG3 #( .INIT(8'h27) )  \bitalign_curr_state_34_4_0_.m23_1_2  (.A(
        late_last_set15_Z), .B(late_flags_pmux), .C(N_20), .Y(m23_1_2));
    CFG4 #( .INIT(16'h2000) )  bitalign_curr_state162 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state161_2_Z), .D(bitalign_curr_state_Z[0]), .Y(
        bitalign_curr_state162_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[105]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[105]), .C(
        un10_early_flags[105]), .Y(early_flags_7_fast_Z[105]));
    SLE \late_flags[5]  (.D(late_flags_7_fast_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[104]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[104]), .C(
        un10_early_flags[104]), .Y(early_flags_7_fast_Z[104]));
    SLE \early_flags[91]  (.D(early_flags_7_fast_Z[91]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[91]));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[4]  (.A(
        tapcnt_final_13_Z[5]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[4]), .Y(tapcnt_final_13_1_Z[4]));
    SLE \late_flags[26]  (.D(late_flags_7_fast_Z[26]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[26]));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[4]  (.A(
        no_early_no_late_val_end1_Z[4]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[4]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[4]));
    ARI1 #( .INIT(20'h51045) )  tapcnt_final_upd_8_cry_3_0 (.A(
        tap_cnt_Z[3]), .B(mv_dn_fg_0_sqmuxa_i_o2_Z), .C(mv_up_fg_Z), 
        .D(N_100), .FCI(tapcnt_final_upd_8_cry_2), .S(
        tapcnt_final_upd_8[3]), .Y(tapcnt_final_upd_8_cry_3_0_Y), .FCO(
        tapcnt_final_upd_8_cry_3));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[48]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[48]), .C(
        un10_early_flags[48]), .Y(early_flags_7_fast_Z[48]));
    CFG3 #( .INIT(8'hF8) )  un1_tap_cnt_0_sqmuxa_1 (.A(
        bitalign_curr_state12_Z), .B(bitalign_curr_state148_Z), .C(
        bitalign_curr_state_1_sqmuxa_4_Z), .Y(un1_tap_cnt_0_sqmuxa_6_0)
        );
    CFG4 #( .INIT(16'h71F9) )  \bitalign_curr_state_34_4_0_.m37_1_1  (
        .A(bitalign_curr_state_Z[1]), .B(bitalign_curr_state_Z[0]), .C(
        early_flags_pmux), .D(N_35), .Y(m37_1_1));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_3 (.A(
        un16_tapcnt_final_3), .B(un10_tapcnt_final_3), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_2_Z), .S(
        un16_tapcnt_final_cry_3_S), .Y(un16_tapcnt_final_cry_3_Y), 
        .FCO(un16_tapcnt_final_cry_3_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_43 (.A(
        un10_early_flags_2_0[40]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_1_Z[40]), .Y(un10_early_flags[43]));
    SLE \wait_cnt[1]  (.D(wait_cnt_4_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(wait_cnt_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[99]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[99]), .C(
        un10_early_flags[99]), .Y(late_flags_7_fast_Z[99]));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[5]  (.A(
        tapcnt_final_13_Z[6]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[5]), .Y(tapcnt_final_13_1_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[45]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[45]), .C(
        un10_early_flags[45]), .Y(early_flags_7_fast_Z[45]));
    CFG4 #( .INIT(16'h4000) )  un10_early_flags_89 (.A(tap_cnt_Z[5]), 
        .B(un10_early_flags_1_Z[9]), .C(un10_early_flags_1_Z[80]), .D(
        un10_early_flags_2_Z[8]), .Y(un10_early_flags[89]));
    CFG2 #( .INIT(4'h2) )  tapcnt_final_upd_2_sqmuxa_1_0_a2_RNO (.A(
        N_100), .B(mv_up_fg_Z), .Y(tapcnt_final_upd_1_sqmuxa));
    ARI1 #( .INIT(20'h45500) )  noearly_nolate_diff_nxt_8_s_7 (.A(VCC), 
        .B(un1_restart_trng_fg_5_Z), .C(GND), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_6), .S(
        noearly_nolate_diff_nxt_8[7]), .Y(
        noearly_nolate_diff_nxt_8_s_7_Y), .FCO(
        noearly_nolate_diff_nxt_8_s_7_FCO));
    CFG4 #( .INIT(16'hFEFF) )  un1_bitalign_curr_state_12 (.A(
        early_flags_1_sqmuxa_1_Z), .B(early_flags_0_sqmuxa_1_Z), .C(
        bitalign_curr_state_Z[1]), .D(un1_bitalign_curr_state148_3_Z), 
        .Y(un1_bitalign_curr_state_12_Z));
    CFG3 #( .INIT(8'hFE) )  un1_bitalign_curr_state_0_sqmuxa_9 (.A(
        rx_err_1_sqmuxa_Z), .B(calc_done_4_sqmuxa_0_Z), .C(
        un1_bitalign_curr_state_0_sqmuxa_9_4_Z), .Y(
        un1_bitalign_curr_state_0_sqmuxa_9_i));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[118]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[118]), .C(
        un10_early_flags[118]), .Y(early_flags_7_fast_Z[118]));
    CFG4 #( .INIT(16'h1000) )  bitalign_curr_state156 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state152_1_Z), .D(bitalign_curr_state_Z[2]), .Y(
        bitalign_curr_state156_Z));
    CFG4 #( .INIT(16'h0080) )  bitalign_curr_state_0_sqmuxa_8 (.A(
        bitalign_curr_state41_Z), .B(bitalign_curr_state152_3_Z), .C(
        BIT_ALGN_OOR_c), .D(bitalign_curr_state_Z[3]), .Y(
        bitalign_curr_state_0_sqmuxa_8_Z));
    SLE \late_flags[76]  (.D(late_flags_7_fast_Z[76]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[76]));
    CFG2 #( .INIT(4'h2) )  \bitalign_curr_state_34_4_0_.m55_0  (.A(
        bitalign_curr_state161_2_Z), .B(bitalign_curr_state_Z[0]), .Y(
        m55_0));
    CFG2 #( .INIT(4'h2) )  early_late_diff_2_sqmuxa (.A(
        early_late_diff_0_sqmuxa_Z), .B(restart_trng_fg_i), .Y(
        early_late_diff_2_sqmuxa_Z));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_95 (.A(
        un10_early_flags_1_Z[80]), .B(tap_cnt_Z[5]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[95]));
    CFG3 #( .INIT(8'h10) )  \bitalign_curr_state_34_4_0_.m52  (.A(
        late_last_set15_Z), .B(early_flags_dec[127]), .C(N_20), .Y(
        N_119_mux));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[77]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[77]), .C(
        un10_early_flags[77]), .Y(late_flags_7_fast_Z[77]));
    SLE reset_dly_fg (.D(VCC), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(reset_dly_fg4_Z), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(reset_dly_fg_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_1_wmux_0 (.A(
        late_flags_pmux_63_1_1_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[32]), .D(late_flags_Z[96]), .FCI(
        late_flags_pmux_63_1_1_co0), .S(
        late_flags_pmux_63_1_1_wmux_0_S), .Y(late_flags_pmux_63_1_1_y1)
        , .FCO(late_flags_pmux_63_1_1_co1));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[111]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[111]), .C(
        un10_early_flags[111]), .Y(early_flags_7_fast_Z[111]));
    ARI1 #( .INIT(20'h0FA44) )  
        \bitalign_curr_state_34_4_0_.m74_2_1_1_1_wmux  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        N_69), .D(m74_1_0), .FCI(VCC), .S(m74_2_1_1_1_wmux_S), .Y(
        m74_2_1_1_1_y0), .FCO(m74_2_1_1_1_co0));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_8_2 (.A(tap_cnt_Z[1]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[8]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[32]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[32]), .C(
        un10_early_flags[32]), .Y(early_flags_7_fast_Z[32]));
    CFG4 #( .INIT(16'hFFFE) )  un2_early_late_diff_validlto7_2 (.A(
        early_late_diff_Z[7]), .B(early_late_diff_Z[6]), .C(
        early_late_diff_Z[5]), .D(early_late_diff_Z[4]), .Y(
        un2_early_late_diff_validlto7_2_Z));
    ARI1 #( .INIT(20'h0FA0C) )  late_flags_pmux_126_1_1_wmux_8 (.A(
        late_flags_pmux_126_1_1_y0_3), .B(late_flags_pmux_126_1_1_y3), 
        .C(late_flags_pmux_126_1_1_y1), .D(emflag_cnt_Z[3]), .FCI(
        late_flags_pmux_126_1_1_co0_3), .S(
        late_flags_pmux_126_1_1_wmux_8_S), .Y(
        late_flags_pmux_126_1_1_y9), .FCO(
        late_flags_pmux_126_1_1_co1_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[31]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[31]), .C(
        un10_early_flags[31]), .Y(late_flags_7_fast_Z[31]));
    SLE \late_flags[7]  (.D(late_flags_7_fast_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[7]));
    CFG4 #( .INIT(16'h0400) )  \bitalign_curr_state_34_4_0_.m91_2  (.A(
        bitalign_curr_state_Z[1]), .B(tap_cnt_0_sqmuxa_0_Z), .C(
        calc_done_Z), .D(bitalign_curr_state_Z[2]), .Y(m91_1));
    CFG4 #( .INIT(16'h8000) )  calc_done25_236 (.A(calc_done25_179_Z), 
        .B(calc_done25_178_Z), .C(calc_done25_177_Z), .D(
        calc_done25_176_Z), .Y(calc_done25_236_Z));
    SLE \late_flags[36]  (.D(late_flags_7_fast_Z[36]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[36]));
    SLE \late_flags[57]  (.D(late_flags_7_fast_Z[57]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[57]));
    CFG4 #( .INIT(16'hF2F0) )  un1_early_flags_1_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(mv_dn_fg_Z), .C(
        early_flags_1_sqmuxa_Z), .D(bitalign_curr_state156_Z), .Y(
        un1_early_flags_1_sqmuxa_i));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_32 (.A(
        un10_early_flags_1_Z[32]), .B(un10_early_flags_2_Z[8]), .C(
        un10_early_flags_2_0[32]), .Y(un10_early_flags[32]));
    CFG4 #( .INIT(16'hFEFA) )  rx_err_1_sqmuxa_RNI2JPB1 (.A(
        timeout_cntlde_0), .B(un1_retrain_adj_tap_i), .C(
        rx_err_1_sqmuxa_Z), .D(N_100), .Y(timeout_cnte));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_3 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[11]), 
        .D(late_flags_Z[75]), .FCI(late_flags_pmux_126_1_0_co1_0), .S(
        late_flags_pmux_126_1_0_wmux_3_S), .Y(
        late_flags_pmux_126_1_0_y0_1), .FCO(
        late_flags_pmux_126_1_0_co0_1));
    ARI1 #( .INIT(20'h54411) )  early_late_diff_8_cry_5_0 (.A(
        emflag_cnt_Z[5]), .B(un1_restart_trng_fg_5_Z), .C(
        early_val_Z[5]), .D(GND), .FCI(early_late_diff_8_cry_4), .S(
        early_late_diff_8[5]), .Y(early_late_diff_8_cry_5_0_Y), .FCO(
        early_late_diff_8_cry_5));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[21]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[21]), .C(
        un10_early_flags[21]), .Y(late_flags_7_fast_Z[21]));
    SLE \late_flags[21]  (.D(late_flags_7_fast_Z[21]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[21]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_cry[1]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[1]), .D(GND), .FCI(
        emflag_cnt_cry_Z[0]), .S(emflag_cnt_s[1]), .Y(
        emflag_cnt_cry_Y_0[1]), .FCO(emflag_cnt_cry_Z[1]));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_cry_3 (.A(
        un10_tapcnt_final_3), .B(early_late_diff_Z[3]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_cry_2_Z), .S(
        un1_early_late_diff_cry_3_S), .Y(un1_early_late_diff_cry_3_Y), 
        .FCO(un1_early_late_diff_cry_3_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[96]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[96]), .C(
        un10_early_flags[96]), .Y(late_flags_7_fast_Z[96]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[1]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[1]), .C(
        un10_early_flags[1]), .Y(late_flags_7_fast_Z[1]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[96]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[96]), .C(
        un10_early_flags[96]), .Y(early_flags_7_fast_Z[96]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_143 (.A(late_flags_Z[75]), 
        .B(late_flags_Z[74]), .C(late_flags_Z[73]), .D(
        late_flags_Z[72]), .Y(calc_done25_143_Z));
    SLE \tapcnt_final[6]  (.D(tapcnt_final_13_1_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[0]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[0]), .C(
        un10_early_flags[0]), .Y(late_flags_7_fast_Z[0]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_1_wmux_14 (.A(
        late_flags_pmux_126_1_1_y0_5), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[53]), .D(late_flags_Z[117]), .FCI(
        late_flags_pmux_126_1_1_co0_6), .S(
        late_flags_pmux_126_1_1_wmux_14_S), .Y(
        late_flags_pmux_126_1_1_y3_0), .FCO(
        late_flags_pmux_126_1_1_co1_6));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_77 (.A(
        un10_early_flags_2_0[76]), .B(un10_early_flags_1_Z[72]), .C(
        un10_early_flags_1_Z[5]), .Y(un10_early_flags[77]));
    CFG4 #( .INIT(16'hF400) )  bit_align_done_0_sqmuxa_2 (.A(
        un1_retrain_adj_tap_i), .B(un1_rx_BIT_ALGN_START), .C(
        bitalign_curr_state12_Z), .D(bitalign_curr_state148_Z), .Y(
        bit_align_done_0_sqmuxa_2_Z));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[17]), 
        .D(late_flags_Z[81]), .FCI(late_flags_pmux_126_1_1_co1), .S(
        late_flags_pmux_126_1_1_wmux_1_S), .Y(
        late_flags_pmux_126_1_1_y0_0), .FCO(
        late_flags_pmux_126_1_1_co0_0));
    CFG4 #( .INIT(16'h3C5A) )  bitalign_curr_state61_3 (.A(
        tapcnt_final_upd_Z[3]), .B(tapcnt_final_Z[3]), .C(tap_cnt_Z[3])
        , .D(N_1416), .Y(bitalign_curr_state61_3_Z));
    ARI1 #( .INIT(20'h44400) )  \timeout_cnt_RNI8UO41[1]  (.A(VCC), .B(
        restart_trng_fg_i), .C(timeout_cnt_Z[1]), .D(GND), .FCI(
        timeout_cnt_cry[0]), .S(timeout_cnt_s[1]), .Y(
        timeout_cnt_RNI8UO41_Y[1]), .FCO(timeout_cnt_cry[1]));
    CFG2 #( .INIT(4'h2) )  un10_early_flags_96_2_0 (.A(
        un10_early_flags_2_Z[0]), .B(tap_cnt_Z[4]), .Y(
        un10_early_flags_2_0[96]));
    SLE \early_flags[88]  (.D(early_flags_7_fast_Z[88]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[88]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_169 (.A(early_flags_Z[83]), 
        .B(early_flags_Z[82]), .C(early_flags_Z[81]), .D(
        early_flags_Z[80]), .Y(calc_done25_169_Z));
    SLE \early_late_diff[0]  (.D(early_late_diff_8[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        early_late_diff_Z[0]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_0 (.A(
        un10_tapcnt_final_0), .B(un16_tapcnt_final_0), .C(GND), .D(GND)
        , .FCI(GND), .S(un10_tapcnt_final_cry_0_S), .Y(
        un10_tapcnt_final_cry_0_Y), .FCO(un10_tapcnt_final_cry_0_Z));
    SLE \noearly_nolate_diff_nxt[6]  (.D(noearly_nolate_diff_nxt_8[6]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_6));
    SLE \tapcnt_final[1]  (.D(tapcnt_final_13_1_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[1]));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_126_1_0_wmux_0 (.A(
        late_flags_pmux_126_1_0_0_y0), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[35]), .D(late_flags_Z[99]), .FCI(
        late_flags_pmux_126_1_0_0_co0), .S(
        late_flags_pmux_126_1_0_wmux_0_S), .Y(
        late_flags_pmux_126_1_0_0_y1), .FCO(
        late_flags_pmux_126_1_0_0_co1));
    SLE \cnt[1]  (.D(cnt_RNO_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(cnt_Z[1]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_22 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_2_0[16]), .C(
        un10_early_flags_1_Z[16]), .Y(un10_early_flags[22]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[121]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[121]), .C(
        un10_early_flags[121]), .Y(late_flags_7_fast_Z[121]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[9]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[9]), .C(
        un10_early_flags[9]), .Y(late_flags_7_fast_Z[9]));
    SLE \late_flags[4]  (.D(late_flags_7_fast_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[4]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_start_7_cry_0_0 (
        .A(emflag_cnt_Z[0]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st1_Z[0]), .D(GND), .FCI(
        noearly_nolate_diff_start_7_cry_0_0_cy_Z), .S(
        noearly_nolate_diff_start_7[0]), .Y(
        noearly_nolate_diff_start_7_cry_0_0_Y), .FCO(
        noearly_nolate_diff_start_7_cry_0));
    SLE \late_flags[71]  (.D(late_flags_7_fast_Z[71]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[71]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[7]), 
        .D(early_flags_Z[71]), .FCI(early_flags_pmux_126_1_0_co1_4), 
        .S(early_flags_pmux_126_1_0_wmux_11_S), .Y(
        early_flags_pmux_126_1_0_y0_4), .FCO(
        early_flags_pmux_126_1_0_co0_5));
    CFG3 #( .INIT(8'h1B) )  \bitalign_curr_state_34_4_0_.m82  (.A(
        bitalign_curr_state_Z[0]), .B(m82_1_0), .C(m82_1_1), .Y(N_83));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_2 (.A(
        early_flags_pmux_63_1_0_y0_0), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[50]), .D(early_flags_Z[114]), .FCI(
        early_flags_pmux_63_1_0_co0_0), .S(
        early_flags_pmux_63_1_0_wmux_2_S), .Y(
        early_flags_pmux_63_1_0_0_y3), .FCO(
        early_flags_pmux_63_1_0_co1_0));
    CFG4 #( .INIT(16'h0001) )  calc_done25_183 (.A(early_flags_Z[43]), 
        .B(early_flags_Z[42]), .C(early_flags_Z[41]), .D(
        early_flags_Z[40]), .Y(calc_done25_183_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[27]), 
        .D(early_flags_Z[91]), .FCI(early_flags_pmux_126_1_0_co1_1), 
        .S(early_flags_pmux_126_1_0_wmux_5_S), .Y(
        early_flags_pmux_126_1_0_y0_2), .FCO(
        early_flags_pmux_126_1_0_co0_2));
    SLE \early_flags[1]  (.D(early_flags_7_fast_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[1]));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_0_2 (.A(tap_cnt_Z[3]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_2_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[53]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[53]), .C(
        un10_early_flags[53]), .Y(early_flags_7_fast_Z[53]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[41]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[41]), .C(
        un10_early_flags[41]), .Y(late_flags_7_fast_Z[41]));
    SLE \tapcnt_final[5]  (.D(tapcnt_final_13_1_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(tapcnt_final_Z[5]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_5 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[27]), 
        .D(late_flags_Z[91]), .FCI(late_flags_pmux_126_1_0_co1_1), .S(
        late_flags_pmux_126_1_0_wmux_5_S), .Y(
        late_flags_pmux_126_1_0_y0_2), .FCO(
        late_flags_pmux_126_1_0_co0_2));
    SLE \late_flags[67]  (.D(late_flags_7_fast_Z[67]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[67]));
    SLE \no_early_no_late_val_end2[4]  (.D(emflag_cnt_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end2_Z[4]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_98 (.A(tap_cnt_Z[1]), 
        .B(tap_cnt_Z[5]), .C(un10_early_flags_1_Z[64]), .D(
        un10_early_flags_2_0[96]), .Y(un10_early_flags[98]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_253 (.A(calc_done25_234_Z), 
        .B(calc_done25_235_Z), .C(calc_done25_251_Z), .D(
        calc_done25_244_Z), .Y(calc_done25_253_Z));
    CFG4 #( .INIT(16'h0001) )  calc_done25_133 (.A(late_flags_Z[99]), 
        .B(late_flags_Z[98]), .C(late_flags_Z[97]), .D(
        late_flags_Z[96]), .Y(calc_done25_133_Z));
    CFG3 #( .INIT(8'hEA) )  un2_noearly_nolate_diff_nxt_validlto2 (.A(
        un16_tapcnt_final_2), .B(un16_tapcnt_final_1), .C(
        un16_tapcnt_final_0), .Y(un2_noearly_nolate_diff_nxt_validlt3));
    SLE \restart_reg[0]  (.D(debouncer_0_DB_OUT), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(restart_reg_Z[0]));
    SLE \early_flags[35]  (.D(early_flags_7_fast_Z[35]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[35]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_19 (.A(tap_cnt_Z[4]), 
        .B(tap_cnt_Z[2]), .C(un10_early_flags_1_Z[3]), .D(
        un10_early_flags_2_0[16]), .Y(un10_early_flags[19]));
    CFG4 #( .INIT(16'hCA42) )  \bitalign_curr_state_34_4_0_.m64  (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[1]), .C(
        m64_1_1), .D(N_63), .Y(N_65));
    ARI1 #( .INIT(20'h5AA55) )  un1_early_late_diff_1_cry_5 (.A(
        un16_tapcnt_final_5), .B(early_late_diff_Z[5]), .C(GND), .D(
        GND), .FCI(un1_early_late_diff_1_cry_4_Z), .S(
        un1_early_late_diff_1_cry_5_S), .Y(
        un1_early_late_diff_1_cry_5_Y), .FCO(
        un1_early_late_diff_1_cry_5_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_9 (.A(
        VCC), .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_126_1_1_co1_3), .S(
        early_flags_pmux_126_1_1_wmux_9_S), .Y(
        early_flags_pmux_126_1_1_wmux_9_Y), .FCO(
        early_flags_pmux_126_1_1_co0_4));
    SLE \late_flags[80]  (.D(late_flags_7_fast_Z[80]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[80]));
    CFG2 #( .INIT(4'h2) )  bit_align_dly_done_2_sqmuxa (.A(
        bitalign_curr_state_0_sqmuxa_9_Z), .B(restart_trng_fg_i), .Y(
        bit_align_dly_done_2_sqmuxa_Z));
    SLE \late_flags[31]  (.D(late_flags_7_fast_Z[31]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[31]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[117]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[117]), .C(
        un10_early_flags[117]), .Y(early_flags_7_fast_Z[117]));
    SLE \early_flags[98]  (.D(early_flags_7_fast_Z[98]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[98]));
    CFG4 #( .INIT(16'h0421) )  un1_bitalign_curr_state148_3 (.A(
        bitalign_curr_state_Z[4]), .B(bitalign_curr_state_Z[3]), .C(
        bitalign_curr_state_Z[0]), .D(bitalign_curr_state_Z[2]), .Y(
        un1_bitalign_curr_state148_3_Z));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_76 (.A(
        un10_early_flags_1_Z[64]), .B(un10_early_flags_2_0[76]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[76]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_115 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[3]), .D(un10_early_flags_2_Z[67]), .Y(
        un10_early_flags[115]));
    SLE \no_early_no_late_val_st1[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_st1_0_sqmuxa_i_Z), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_st1_Z[0]));
    CFG4 #( .INIT(16'hFFF1) )  un1_bitalign_curr_state148_8_2 (.A(
        un1_bitalign_curr_state148_5_4_Z), .B(
        un1_bitalign_curr_state148_4_1_Z), .C(
        un1_bitalign_curr_state148_8_0_Z), .D(rx_trng_done_1_sqmuxa_Z), 
        .Y(un1_bitalign_curr_state148_8_2_Z));
    ARI1 #( .INIT(20'h0F588) )  late_flags_pmux_63_1_0_wmux_4 (.A(
        late_flags_pmux_63_1_0_y0_1), .B(emflag_cnt_Z[5]), .C(
        late_flags_Z[42]), .D(late_flags_Z[106]), .FCI(
        late_flags_pmux_63_1_0_co0_1), .S(
        late_flags_pmux_63_1_0_wmux_4_S), .Y(
        late_flags_pmux_63_1_0_0_y5), .FCO(
        late_flags_pmux_63_1_0_co1_1));
    SLE \rst_cnt[5]  (.D(rst_cnt_s[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[5]));
    CFG4 #( .INIT(16'hFF8C) )  un1_restart_trng_fg_10 (.A(
        calc_done25_Z), .B(bitalign_curr_state162_Z), .C(
        un1_calc_done25_7_i), .D(un1_restart_trng_fg_10_0_Z), .Y(
        un1_restart_trng_fg_10_sn));
    SLE \tap_cnt[0]  (.D(N_32_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G)
        , .EN(VCC), .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), 
        .SD(GND), .LAT(GND), .Q(tap_cnt_Z[0]));
    SLE \no_early_no_late_val_end1[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[0]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[33]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[33]), .C(
        un10_early_flags[33]), .Y(late_flags_7_fast_Z[33]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[43]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[43]), .C(
        un10_early_flags[43]), .Y(early_flags_7_fast_Z[43]));
    SLE \late_flags[10]  (.D(late_flags_7_fast_Z[10]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[10]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[102]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[102]), .C(
        un10_early_flags[102]), .Y(early_flags_7_fast_Z[102]));
    ARI1 #( .INIT(20'h5AA55) )  un10_tapcnt_final_cry_7 (.A(
        un10_tapcnt_final_7), .B(un16_tapcnt_final_7), .C(GND), .D(GND)
        , .FCI(un10_tapcnt_final_cry_6_Z), .S(
        un10_tapcnt_final_cry_7_S), .Y(un10_tapcnt_final_cry_7_Y), 
        .FCO(un10_tapcnt_final_cry_7_Z));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNID5OPG[4]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNIPMIR_Z[4]), .B(
        early_val_RNIF13D1_Z[4]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[4]), .FCI(tapcnt_final_13_m1_cry_3), .S(
        tapcnt_final_13_m1[4]), .Y(early_val_RNID5OPG_Y[4]), .FCO(
        tapcnt_final_13_m1_cry_4));
    CFG2 #( .INIT(4'h8) )  un10_early_flags_6_1 (.A(tap_cnt_Z[1]), .B(
        tap_cnt_Z[2]), .Y(un10_early_flags_1_Z[6]));
    SLE \early_flags[65]  (.D(early_flags_7_fast_Z[65]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[65]));
    CFG2 #( .INIT(4'h2) )  \tap_cnt_RNO[3]  (.A(N_77), .B(N_63_0), .Y(
        N_26_i));
    ARI1 #( .INIT(20'h572D8) )  \tapcnt_final_RNI2SF33[2]  (.A(
        un1_tap_cnt_0_sqmuxa_14_0_Z[1]), .B(N_60), .C(tap_cnt_Z[2]), 
        .D(tapcnt_final_Z[2]), .FCI(tap_cnt_17_i_m2_cry_1), .S(N_78), 
        .Y(tapcnt_final_RNI2SF33_Y[2]), .FCO(tap_cnt_17_i_m2_cry_2));
    SLE \bitalign_curr_state[2]  (.D(bitalign_curr_state_34[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(bitalign_curr_state_Z[2]));
    ARI1 #( .INIT(20'h574B8) )  \tapcnt_final_RNIES844[3]  (.A(
        tap_cnt_Z[3]), .B(un1_tap_cnt_0_sqmuxa_14_0_Z[1]), .C(N_60), 
        .D(tapcnt_final_Z[3]), .FCI(tap_cnt_17_i_m2_cry_2), .S(N_77), 
        .Y(tapcnt_final_RNIES844_Y[3]), .FCO(tap_cnt_17_i_m2_cry_3));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[23]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[23]), .C(
        un10_early_flags[23]), .Y(late_flags_7_fast_Z[23]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_174 (.A(early_flags_Z[79]), 
        .B(early_flags_Z[78]), .C(early_flags_Z[77]), .D(
        early_flags_Z[76]), .Y(calc_done25_174_Z));
    SLE \late_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[6])
        );
    SLE \early_val[6]  (.D(emflag_cnt_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_val_0_sqmuxa_1_i_Z)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_val_Z[6]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[21]), 
        .D(early_flags_Z[85]), .FCI(early_flags_pmux_126_1_1_co1_5), 
        .S(early_flags_pmux_126_1_1_wmux_13_S), .Y(
        early_flags_pmux_126_1_1_y0_5), .FCO(
        early_flags_pmux_126_1_1_co0_6));
    SLE \tapcnt_final_upd[0]  (.D(tapcnt_final_upd_8_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[0]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_0_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[7]), .D(
        late_flags_Z[71]), .FCI(late_flags_pmux_126_1_0_co1_4), .S(
        late_flags_pmux_126_1_0_wmux_11_S), .Y(
        late_flags_pmux_126_1_0_y0_4), .FCO(
        late_flags_pmux_126_1_0_co0_5));
    SLE \late_flags[40]  (.D(late_flags_7_fast_Z[40]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[40]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[30]), 
        .D(late_flags_Z[94]), .FCI(late_flags_pmux_63_1_0_co1_7), .S(
        late_flags_pmux_63_1_0_wmux_17_S), .Y(
        late_flags_pmux_63_1_0_y0_7), .FCO(
        late_flags_pmux_63_1_0_co0_8));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_91 (.A(
        un10_early_flags_1_Z[24]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[5]), .D(un10_early_flags_2_Z[67]), .Y(
        un10_early_flags[91]));
    CFG4 #( .INIT(16'hFFFE) )  un34lto7_4 (.A(un16_tapcnt_final_3), .B(
        un16_tapcnt_final_2), .C(un16_tapcnt_final_1), .D(
        un16_tapcnt_final_0), .Y(un34lto7_4_Z));
    CFG2 #( .INIT(4'h2) )  rx_BIT_ALGN_DIR_1_sqmuxa (.A(
        bitalign_curr_state155_Z), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(rx_BIT_ALGN_DIR_1_sqmuxa_Z));
    SLE \early_flags[108]  (.D(early_flags_7_fast_Z[108]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[108]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_35 (.A(
        un10_early_flags_2_0[32]), .B(un10_early_flags_1_Z[3]), .C(
        un10_early_flags_2_Z[35]), .Y(un10_early_flags[35]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[70]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[70]), .C(
        un10_early_flags[70]), .Y(late_flags_7_fast_Z[70]));
    SLE \late_flags[116]  (.D(late_flags_7_fast_Z[116]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[116]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[9]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[9]), .C(
        un10_early_flags[9]), .Y(early_flags_7_fast_Z[9]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_53 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[5]), .C(
        un10_early_flags_2_0[52]), .Y(un10_early_flags[53]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_149 (.A(late_flags_Z[35]), 
        .B(late_flags_Z[34]), .C(late_flags_Z[33]), .D(
        late_flags_Z[32]), .Y(calc_done25_149_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[37]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[37]), .C(
        un10_early_flags[37]), .Y(early_flags_7_fast_Z[37]));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_105 (.A(
        un10_early_flags_1_Z[9]), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[96]), .D(un10_early_flags_2_Z[8]), .Y(
        un10_early_flags[105]));
    CFG4 #( .INIT(16'h0400) )  bitalign_curr_state_1_sqmuxa_7_0_a2_0 (
        .A(bitalign_curr_state12_Z), .B(bitalign_curr_state148_Z), .C(
        BIT_ALGN_ERR_0_c), .D(retrain_reg_Z[2]), .Y(N_100));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_1_wmux_6 (.A(
        early_flags_pmux_63_1_1_y0_2), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[56]), .D(early_flags_Z[120]), .FCI(
        early_flags_pmux_63_1_1_co0_2), .S(
        early_flags_pmux_63_1_1_wmux_6_S), .Y(
        early_flags_pmux_63_1_1_y7), .FCO(
        early_flags_pmux_63_1_1_co1_2));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_11 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[5]), .D(
        late_flags_Z[69]), .FCI(late_flags_pmux_126_1_1_co1_4), .S(
        late_flags_pmux_126_1_1_wmux_11_S), .Y(
        late_flags_pmux_126_1_1_y0_4), .FCO(
        late_flags_pmux_126_1_1_co0_5));
    SLE \late_val[0]  (.D(emflag_cnt_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        early_late_diff_0_sqmuxa_1_i), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(N_19_i), .SD(GND), .LAT(GND), .Q(late_val_Z[0])
        );
    CFG3 #( .INIT(8'h74) )  un1_bitalign_curr_state152 (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[0]), .C(
        bitalign_curr_state155_1_Z), .Y(un1_bitalign_curr_state152_Z));
    SLE \tapcnt_final_upd[6]  (.D(tapcnt_final_upd_8[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        tapcnt_final_upd_0_sqmuxa_i_Z), .ALn(RX_CLK_ALIGN_DONE_arst), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        tapcnt_final_upd_Z[6]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[43]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[43]), .C(
        un10_early_flags[43]), .Y(late_flags_7_fast_Z[43]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_126_1_1_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[17]), 
        .D(early_flags_Z[81]), .FCI(early_flags_pmux_126_1_1_co1), .S(
        early_flags_pmux_126_1_1_wmux_1_S), .Y(
        early_flags_pmux_126_1_1_y0_0), .FCO(
        early_flags_pmux_126_1_1_co0_0));
    CFG4 #( .INIT(16'hC505) )  \bitalign_curr_state_34_4_0_.m10  (.A(
        BIT_ALGN_OOR_c), .B(calc_done_Z), .C(bitalign_curr_state_Z[0]), 
        .D(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .Y(N_11));
    SLE \no_early_no_late_val_st2[1]  (.D(emflag_cnt_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(un1_restart_trng_fg_8_Z), 
        .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND)
        , .LAT(GND), .Q(no_early_no_late_val_st2_Z[1]));
    CFG3 #( .INIT(8'h1D) )  \no_early_no_late_val_st1_RNIV8921[3]  (.A(
        no_early_no_late_val_st1_Z[3]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_st2_Z[3]), .Y(
        un1_no_early_no_late_val_st1_1_1[3]));
    SLE \noearly_nolate_diff_nxt[3]  (.D(noearly_nolate_diff_nxt_8[3]), 
        .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end2_0_sqmuxa_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un16_tapcnt_final_3));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNINKIR[3]  (.A(
        late_val_Z[3]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[3]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNINKIR_Z[3]));
    SLE \early_flags[6]  (.D(early_flags_7_fast_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[6]));
    CFG4 #( .INIT(16'h0800) )  un10_early_flags_63 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[63]));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNILIIR[2]  (.A(
        late_val_Z[2]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[2]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNILIIR_Z[2]));
    SLE \early_flags[75]  (.D(early_flags_7_fast_Z[75]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[75]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_25 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_0[24]), .C(
        un10_early_flags_2_Z[21]), .Y(un10_early_flags[25]));
    SLE \early_flags[53]  (.D(early_flags_7_fast_Z[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[53]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_189 (.A(early_flags_Z[3]), 
        .B(early_flags_Z[2]), .C(early_flags_Z[1]), .D(
        early_flags_Z[0]), .Y(calc_done25_189_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[108]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[108]), .C(
        un10_early_flags[108]), .Y(early_flags_7_fast_Z[108]));
    CFG4 #( .INIT(16'hFFFE) )  
        un2_noearly_nolate_diff_start_validlto7_2 (.A(
        un10_tapcnt_final_7), .B(un10_tapcnt_final_6), .C(
        un10_tapcnt_final_5), .D(un10_tapcnt_final_4), .Y(
        un2_noearly_nolate_diff_start_validlto7_2_Z));
    CFG3 #( .INIT(8'h8B) )  
        \un1_no_early_no_late_val_end1_1_1_RNIPMIR[4]  (.A(
        late_val_Z[4]), .B(tapcnt_final_3_sqmuxa_Z), .C(
        un1_no_early_no_late_val_end1_1_1_Z[4]), .Y(
        un1_no_early_no_late_val_end1_1_1_RNIPMIR_Z[4]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_139 (.A(late_flags_Z[91]), 
        .B(late_flags_Z[90]), .C(late_flags_Z[89]), .D(
        late_flags_Z[88]), .Y(calc_done25_139_Z));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[20]), 
        .D(early_flags_Z[84]), .FCI(early_flags_pmux_63_1_1_co1_5), .S(
        early_flags_pmux_63_1_1_wmux_13_S), .Y(
        early_flags_pmux_63_1_1_y0_5), .FCO(
        early_flags_pmux_63_1_1_co0_6));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[76]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[76]), .C(
        un10_early_flags[76]), .Y(early_flags_7_fast_Z[76]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[101]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[101]), .C(
        un10_early_flags[101]), .Y(early_flags_7_fast_Z[101]));
    CFG3 #( .INIT(8'hE4) )  \late_flags_RNO[49]  (.A(N_208), .B(
        EYE_MONITOR_LATE_net_0_0), .C(late_flags_Z[49]), .Y(
        late_flags_RNO_Z[49]));
    ARI1 #( .INIT(20'h0FA0C) )  early_flags_pmux_63_1_1_wmux_20 (.A(
        early_flags_pmux_63_1_1_y0_8), .B(early_flags_pmux_63_1_1_y3_0)
        , .C(early_flags_pmux_63_1_1_y1_0), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co0_9), .S(
        early_flags_pmux_63_1_1_wmux_20_S), .Y(
        early_flags_pmux_63_1_1_y21), .FCO(
        early_flags_pmux_63_1_1_co1_9));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_63_1_0_wmux_16 (.A(
        early_flags_pmux_63_1_0_y0_6), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[46]), .D(early_flags_Z[110]), .FCI(
        early_flags_pmux_63_1_0_co0_7), .S(
        early_flags_pmux_63_1_0_wmux_16_S), .Y(
        early_flags_pmux_63_1_0_y5_0), .FCO(
        early_flags_pmux_63_1_0_co1_7));
    SLE \early_flags[109]  (.D(early_flags_7_fast_Z[109]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[109]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_9 (.A(
        un10_early_flags_1_Z[9]), .B(un10_early_flags_2_Z[8]), .C(
        un10_early_flags_2_0[0]), .Y(un10_early_flags[9]));
    SLE \noearly_nolate_diff_start[6]  (.D(
        noearly_nolate_diff_start_7[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_6));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[22]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[22]), .C(
        un10_early_flags[22]), .Y(early_flags_7_fast_Z[22]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[58]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[58]), .C(
        un10_early_flags[58]), .Y(late_flags_7_fast_Z[58]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_9 (.A(VCC)
        , .B(VCC), .C(emflag_cnt_Z[2]), .D(VCC), .FCI(
        early_flags_pmux_63_1_1_co1_3), .S(
        early_flags_pmux_63_1_1_wmux_9_S), .Y(
        early_flags_pmux_63_1_1_wmux_9_Y), .FCO(
        early_flags_pmux_63_1_1_co0_4));
    CFG4 #( .INIT(16'h2000) )  un10_early_flags_90 (.A(
        un10_early_flags_1_Z[10]), .B(tap_cnt_Z[5]), .C(
        un10_early_flags_1_Z[80]), .D(un10_early_flags_2_Z[10]), .Y(
        un10_early_flags[90]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[82]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[82]), .C(
        un10_early_flags[82]), .Y(early_flags_7_fast_Z[82]));
    SLE \noearly_nolate_diff_start[2]  (.D(
        noearly_nolate_diff_start_7[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(un10_tapcnt_final_2));
    SLE \early_flags[19]  (.D(early_flags_7_fast_Z[19]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[19]));
    SLE \late_flags[53]  (.D(late_flags_7_fast_Z[53]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[53]));
    SLE \early_flags[20]  (.D(early_flags_7_fast_Z[20]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[20]));
    CFG4 #( .INIT(16'hF6FF) )  un1_bitalign_curr_state_14_1 (.A(
        bitalign_curr_state_Z[2]), .B(bitalign_curr_state_Z[3]), .C(
        tapcnt_final_upd_3_sqmuxa_Z), .D(N_117_mux_1), .Y(
        un1_bitalign_curr_state_14_1_Z));
    SLE \late_flags[90]  (.D(late_flags_7_fast_Z[90]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[90]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[12]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[12]), .C(
        un10_early_flags[12]), .Y(late_flags_7_fast_Z[12]));
    CFG4 #( .INIT(16'h8000) )  calc_done25_227 (.A(calc_done25_143_Z), 
        .B(calc_done25_142_Z), .C(calc_done25_141_Z), .D(
        calc_done25_140_Z), .Y(calc_done25_227_Z));
    CFG4 #( .INIT(16'h8000) )  calc_done25_228 (.A(calc_done25_147_Z), 
        .B(calc_done25_146_Z), .C(calc_done25_145_Z), .D(
        calc_done25_144_Z), .Y(calc_done25_228_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[62]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[62]), .C(
        un10_early_flags[62]), .Y(early_flags_7_fast_Z[62]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_38 (.A(
        un10_early_flags_1_Z[6]), .B(un10_early_flags_2_0[32]), .C(
        un10_early_flags_1_Z[32]), .Y(un10_early_flags[38]));
    ARI1 #( .INIT(20'h574B8) )  \early_val_RNIO46ED[3]  (.A(
        un1_no_early_no_late_val_end1_1_1_RNINKIR_Z[3]), .B(
        early_val_RNICU2D1_Z[3]), .C(un1_bitalign_curr_state169_12_sn), 
        .D(early_val_Z[3]), .FCI(tapcnt_final_13_m1_cry_2), .S(
        tapcnt_final_13_m1[3]), .Y(early_val_RNIO46ED_Y[3]), .FCO(
        tapcnt_final_13_m1_cry_3));
    SLE \late_flags[85]  (.D(late_flags_7_fast_Z[85]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[85]));
    ARI1 #( .INIT(20'h4AA00) )  \rst_cnt_cry[3]  (.A(VCC), .B(
        rst_cnt_Z[3]), .C(GND), .D(GND), .FCI(rst_cnt_cry_Z[2]), .S(
        rst_cnt_s[3]), .Y(rst_cnt_cry_Y_0[3]), .FCO(rst_cnt_cry_Z[3]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[39]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[39]), .C(
        un10_early_flags[39]), .Y(late_flags_7_fast_Z[39]));
    SLE \early_flags[114]  (.D(early_flags_7_fast_Z[114]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[114]));
    CFG3 #( .INIT(8'h5D) )  un1_early_flags_pmux_1_RNIV4F8 (.A(
        early_late_diff_0_sqmuxa_1_0_Z), .B(bitalign_curr_state159_Z), 
        .C(un1_early_flags_pmux_1_Z), .Y(
        no_early_no_late_val_end1_0_sqmuxa_1_i));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_1 (.A(late_val_Z[1])
        , .B(early_val_Z[1]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_0_Z), .S(tapcnt_final27_cry_1_S), .Y(
        tapcnt_final27_cry_1_Y), .FCO(tapcnt_final27_cry_1_Z));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_126_1_1_wmux_7 (.A(
        early_flags_pmux_126_1_1_y7), .B(early_flags_pmux_126_1_1_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_126_1_1_co1_2), .S(
        early_flags_pmux_126_1_1_wmux_7_S), .Y(
        early_flags_pmux_126_1_1_y0_3), .FCO(
        early_flags_pmux_126_1_1_co0_3));
    CFG2 #( .INIT(4'h8) )  tap_cnt_0_sqmuxa_0 (.A(
        bitalign_curr_state_Z[0]), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), 
        .Y(tap_cnt_0_sqmuxa_0_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[8]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[8]), .C(
        un10_early_flags[8]), .Y(late_flags_7_fast_Z[8]));
    CFG4 #( .INIT(16'hA888) )  un2_early_late_diff_validlto3 (.A(
        early_late_diff_Z[3]), .B(early_late_diff_Z[2]), .C(
        early_late_diff_Z[1]), .D(early_late_diff_Z[0]), .Y(
        un2_early_late_diff_validlt7));
    ARI1 #( .INIT(20'h5AA55) )  un16_tapcnt_final_cry_5 (.A(
        un16_tapcnt_final_5), .B(un10_tapcnt_final_5), .C(GND), .D(GND)
        , .FCI(un16_tapcnt_final_cry_4_Z), .S(
        un16_tapcnt_final_cry_5_S), .Y(un16_tapcnt_final_cry_5_Y), 
        .FCO(un16_tapcnt_final_cry_5_Z));
    SLE \rst_cnt[9]  (.D(rst_cnt_s_Z[9]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(rst_cnt_Z[9]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[29]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[29]), .C(
        un10_early_flags[29]), .Y(late_flags_7_fast_Z[29]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[39]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[39]), .C(
        un10_early_flags[39]), .Y(early_flags_7_fast_Z[39]));
    CFG4 #( .INIT(16'hFFFE) )  un1_calc_done25_5 (.A(
        un1_tapcnt_final_Z), .B(un1_noearly_nolate_diff_nxt_valid_Z), 
        .C(calc_done25_Z), .D(un1_noearly_nolate_diff_start_valid_Z), 
        .Y(un1_calc_done25_5_Z));
    SLE \late_flags[15]  (.D(late_flags_7_fast_Z[15]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[15]));
    SLE \early_flags[101]  (.D(early_flags_7_fast_Z[101]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[101]));
    SLE \late_flags[63]  (.D(late_flags_7_fast_Z[63]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[63]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_28 (.A(
        un10_early_flags_2_0[28]), .B(un10_early_flags_1_Z[16]), .C(
        un10_early_flags_1_Z[12]), .Y(un10_early_flags[28]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[10]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[10]), .C(
        un10_early_flags[10]), .Y(early_flags_7_fast_Z[10]));
    CFG4 #( .INIT(16'hFF40) )  un1_rx_BIT_ALGN_LOAD_0_sqmuxa (.A(
        calc_done_Z), .B(sig_rx_BIT_ALGN_CLR_FLGS14_Z), .C(
        bitalign_curr_state154_Z), .D(rx_BIT_ALGN_LOAD_0_sqmuxa_Z), .Y(
        un1_rx_BIT_ALGN_LOAD_0_sqmuxa_i_0));
    CFG3 #( .INIT(8'h20) )  \bitalign_curr_state_34_4_0_.m72  (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state_Z[0]), 
        .C(bitalign_curr_state61), .Y(N_116_mux));
    SLE \early_flags[22]  (.D(early_flags_7_fast_Z[22]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[22]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[78]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[78]), .C(
        un10_early_flags[78]), .Y(late_flags_7_fast_Z[78]));
    CFG2 #( .INIT(4'hE) )  un1_calc_done25_7 (.A(un1_calc_done25_5_Z), 
        .B(un1_early_late_diff_valid_Z), .Y(un1_calc_done25_7_i));
    CFG3 #( .INIT(8'hE2) )  \tapcnt_final_13_1[1]  (.A(
        tapcnt_final_13_Z[2]), .B(un1_tapcnt_final_0_sqmuxa_Z), .C(
        tapcnt_final_13_Z[1]), .Y(tapcnt_final_13_1_Z[1]));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[0]), 
        .D(early_flags_Z[64]), .FCI(VCC), .S(
        early_flags_pmux_63_1_1_wmux_S), .Y(early_flags_pmux_63_1_1_y0)
        , .FCO(early_flags_pmux_63_1_1_co0));
    SLE \early_flags[103]  (.D(early_flags_7_fast_Z[103]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[103]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_127 (.A(
        un10_early_flags_1_Z[48]), .B(un10_early_flags_1_Z[3]), .C(
        tap_cnt_Z[6]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[127]));
    SLE \late_flags[124]  (.D(late_flags_7_fast_Z[124]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[124]));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_4 (.A(late_val_Z[4])
        , .B(early_val_Z[4]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_3_Z), .S(tapcnt_final27_cry_4_S), .Y(
        tapcnt_final27_cry_4_Y), .FCO(tapcnt_final27_cry_4_Z));
    ARI1 #( .INIT(20'h45500) )  restart_trng_fg_RNIBNT7 (.A(VCC), .B(
        restart_trng_fg_i), .C(GND), .D(GND), .FCI(VCC), .S(
        restart_trng_fg_RNIBNT7_S), .Y(restart_trng_fg_RNIBNT7_Y), 
        .FCO(timeout_cnt_cry_cy));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_126_1_1_wmux_13 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[21]), 
        .D(late_flags_Z[85]), .FCI(late_flags_pmux_126_1_1_co1_5), .S(
        late_flags_pmux_126_1_1_wmux_13_S), .Y(
        late_flags_pmux_126_1_1_y0_5), .FCO(
        late_flags_pmux_126_1_1_co0_6));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[112]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[112]), .C(
        un10_early_flags[112]), .Y(late_flags_7_fast_Z[112]));
    SLE \late_flags[45]  (.D(late_flags_7_fast_Z[45]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[45]));
    CFG3 #( .INIT(8'h80) )  sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa (.A(
        sig_rx_BIT_ALGN_CLR_FLGS14_Z), .B(bitalign_curr_state154_Z), 
        .C(calc_done_Z), .Y(sig_rx_BIT_ALGN_CLR_FLGS_0_sqmuxa_Z));
    SLE \late_flags[28]  (.D(late_flags_7_fast_Z[28]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[28]));
    CFG4 #( .INIT(16'h0001) )  calc_done25_160 (.A(early_flags_Z[119]), 
        .B(early_flags_Z[118]), .C(early_flags_Z[117]), .D(
        early_flags_Z[116]), .Y(calc_done25_160_Z));
    CFG4 #( .INIT(16'h0001) )  \un1_tap_cnt_0_sqmuxa_14_i_a2[0]  (.A(
        un1_early_flags_1_sqmuxa_i), .B(rx_BIT_ALGN_MOVE_0_sqmuxa_1_Z), 
        .C(N_63_0), .D(bitalign_curr_state_0_sqmuxa_10), .Y(N_89));
    ARI1 #( .INIT(20'h5AA55) )  tapcnt_final27_cry_3 (.A(late_val_Z[3])
        , .B(early_val_Z[3]), .C(GND), .D(GND), .FCI(
        tapcnt_final27_cry_2_Z), .S(tapcnt_final27_cry_3_S), .Y(
        tapcnt_final27_cry_3_Y), .FCO(tapcnt_final27_cry_3_Z));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[36]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[36]), .C(
        un10_early_flags[36]), .Y(late_flags_7_fast_Z[36]));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[107]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[107]), .C(
        un10_early_flags[107]), .Y(early_flags_7_fast_Z[107]));
    ARI1 #( .INIT(20'h51045) )  tapcnt_final_upd_8_cry_5_0 (.A(
        tap_cnt_Z[5]), .B(mv_dn_fg_0_sqmuxa_i_o2_Z), .C(mv_up_fg_Z), 
        .D(N_100), .FCI(tapcnt_final_upd_8_cry_4), .S(
        tapcnt_final_upd_8[5]), .Y(tapcnt_final_upd_8_cry_5_0_Y), .FCO(
        tapcnt_final_upd_8_cry_5));
    CFG4 #( .INIT(16'h202F) )  \tapcnt_final_13_1_1_0[0]  (.A(
        tapcnt_final_Z[0]), .B(un1_restart_trng_fg_10_sn), .C(
        tapcnt_final_13_m0s2_Z), .D(early_val_RNIT7HB3_Y[0]), .Y(
        tapcnt_final_13_1_1_0_Z[0]));
    CFG2 #( .INIT(4'h2) )  rx_BIT_ALGN_MOVE_2_sqmuxa (.A(
        un1_early_flags_1_sqmuxa_1_Z), .B(restart_trng_fg_i), .Y(
        rx_BIT_ALGN_MOVE_2_sqmuxa_Z));
    SLE \early_flags[83]  (.D(early_flags_7_fast_Z[83]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(early_flags_Z[83]));
    CFG4 #( .INIT(16'h8000) )  un10_early_flags_31 (.A(
        un10_early_flags_30_0_Z), .B(tap_cnt_Z[4]), .C(
        un10_early_flags_1_Z[3]), .D(un10_early_flags_1_Z[12]), .Y(
        un10_early_flags[31]));
    CFG3 #( .INIT(8'h1D) )  \un1_no_early_no_late_val_end1_1_1[5]  (.A(
        no_early_no_late_val_end1_Z[5]), .B(tapcnt_final_2_sqmuxa_Z), 
        .C(no_early_no_late_val_end2_Z[5]), .Y(
        un1_no_early_no_late_val_end1_1_1_Z[5]));
    CFG3 #( .INIT(8'hAC) )  \late_flags_7_fast[26]  (.A(
        EYE_MONITOR_LATE_net_0_0), .B(late_flags_Z[26]), .C(
        un10_early_flags[26]), .Y(late_flags_7_fast_Z[26]));
    ARI1 #( .INIT(20'h48800) )  \emflag_cnt_s[6]  (.A(VCC), .B(
        emflag_cnt_cry_cy_Y_0[0]), .C(emflag_cnt_Z[6]), .D(GND), .FCI(
        emflag_cnt_cry_Z[5]), .S(emflag_cnt_s_Z[6]), .Y(
        emflag_cnt_s_Y[6]), .FCO(emflag_cnt_s_FCO[6]));
    SLE \late_flags[118]  (.D(late_flags_7_fast_Z[118]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[118]));
    ARI1 #( .INIT(20'h0EC2C) )  early_flags_pmux_63_1_1_wmux_7 (.A(
        early_flags_pmux_63_1_1_y7), .B(early_flags_pmux_63_1_1_y5), 
        .C(emflag_cnt_Z[4]), .D(emflag_cnt_Z[3]), .FCI(
        early_flags_pmux_63_1_1_co1_2), .S(
        early_flags_pmux_63_1_1_wmux_7_S), .Y(
        early_flags_pmux_63_1_1_y0_3), .FCO(
        early_flags_pmux_63_1_1_co0_3));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_63_1_1_wmux_17 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(early_flags_Z[28]), 
        .D(early_flags_Z[92]), .FCI(early_flags_pmux_63_1_1_co1_7), .S(
        early_flags_pmux_63_1_1_wmux_17_S), .Y(
        early_flags_pmux_63_1_1_y0_7), .FCO(
        early_flags_pmux_63_1_1_co0_8));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[126]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[126]), .C(
        un10_early_flags[126]), .Y(early_flags_7_fast_Z[126]));
    ARI1 #( .INIT(20'h54411) )  noearly_nolate_diff_nxt_8_cry_6_0 (.A(
        emflag_cnt_Z[6]), .B(un1_restart_trng_fg_5_Z), .C(
        no_early_no_late_val_st2_Z[6]), .D(GND), .FCI(
        noearly_nolate_diff_nxt_8_cry_5), .S(
        noearly_nolate_diff_nxt_8[6]), .Y(
        noearly_nolate_diff_nxt_8_cry_6_0_Y), .FCO(
        noearly_nolate_diff_nxt_8_cry_6));
    ARI1 #( .INIT(20'h0F588) )  early_flags_pmux_126_1_1_wmux_4 (.A(
        early_flags_pmux_126_1_1_y0_1), .B(emflag_cnt_Z[5]), .C(
        early_flags_Z[41]), .D(early_flags_Z[105]), .FCI(
        early_flags_pmux_126_1_1_co0_1), .S(
        early_flags_pmux_126_1_1_wmux_4_S), .Y(
        early_flags_pmux_126_1_1_y5), .FCO(
        early_flags_pmux_126_1_1_co1_1));
    CFG3 #( .INIT(8'h40) )  rx_trng_done_RNO (.A(restart_trng_fg_i), 
        .B(bitalign_curr_state41_Z), .C(bitalign_curr_state_Z[1]), .Y(
        N_1403));
    CFG4 #( .INIT(16'hF1F0) )  rx_trng_done_0_sqmuxa_i (.A(
        early_flags_1_sqmuxa_1_Z), .B(un1_bitalign_curr_state_13_1_Z), 
        .C(restart_trng_fg_i), .D(un1_bitalign_curr_state148_2_Z), .Y(
        rx_trng_done_0_sqmuxa_i_Z));
    SLE \late_flags[78]  (.D(late_flags_7_fast_Z[78]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(early_flags_0_sqmuxa_2_i)
        , .ALn(RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(
        GND), .LAT(GND), .Q(late_flags_Z[78]));
    SLE \no_early_no_late_val_end1[3]  (.D(emflag_cnt_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        no_early_no_late_val_end1_0_sqmuxa_1_i), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(N_19_i), .SD(GND), 
        .LAT(GND), .Q(no_early_no_late_val_end1_Z[3]));
    CFG3 #( .INIT(8'h04) )  bitalign_curr_state155 (.A(
        un1_bitalign_curr_state_15_1_Z), .B(bitalign_curr_state155_1_Z)
        , .C(bitalign_curr_state_Z[3]), .Y(bitalign_curr_state155_Z));
    CFG2 #( .INIT(4'h1) )  un10_early_flags_30_0 (.A(tap_cnt_Z[5]), .B(
        tap_cnt_Z[6]), .Y(un10_early_flags_30_0_Z));
    CFG3 #( .INIT(8'hAC) )  \early_flags_7_fast[14]  (.A(
        EYE_MONITOR_EARLY_net_0_0), .B(early_flags_Z[14]), .C(
        un10_early_flags[14]), .Y(early_flags_7_fast_Z[14]));
    CFG3 #( .INIT(8'h80) )  un10_early_flags_21 (.A(
        un10_early_flags_1_Z[5]), .B(un10_early_flags_2_0[16]), .C(
        un10_early_flags_2_Z[21]), .Y(un10_early_flags[21]));
    ARI1 #( .INIT(20'h0FA44) )  late_flags_pmux_63_1_0_wmux_1 (.A(
        emflag_cnt_Z[6]), .B(emflag_cnt_Z[5]), .C(late_flags_Z[18]), 
        .D(late_flags_Z[82]), .FCI(late_flags_pmux_63_1_0_0_co1), .S(
        late_flags_pmux_63_1_0_wmux_1_S), .Y(
        late_flags_pmux_63_1_0_y0_0), .FCO(
        late_flags_pmux_63_1_0_co0_0));
    ARI1 #( .INIT(20'h0FA44) )  early_flags_pmux_127_1_0_wmux (.A(
        emflag_cnt_Z[1]), .B(emflag_cnt_Z[0]), .C(
        early_flags_pmux_63_1_1_wmux_10_Y), .D(
        early_flags_pmux_63_1_0_wmux_10_Y), .FCI(VCC), .S(
        early_flags_pmux_127_1_0_wmux_S), .Y(
        early_flags_pmux_127_1_0_y0), .FCO(
        early_flags_pmux_127_1_0_co0));
    
endmodule


module 
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_0s_0s_0s_26s_10s_10s_1(
        
       EYE_MONITOR_LATE_net_0_0,
       EYE_MONITOR_EARLY_net_0_0,
       BIT_ALGN_EYE_IN_c,
       RX_CLK_ALIGN_DONE_arst,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       debouncer_0_DB_OUT,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE,
       BIT_ALGN_ERR_0_c,
       BIT_ALGN_OOR_c,
       BIT_ALGN_START_1_c,
       BIT_ALGN_DONE_c,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS,
       PLL_LOCK_0
    );
input  EYE_MONITOR_LATE_net_0_0;
input  EYE_MONITOR_EARLY_net_0_0;
input  [2:0] BIT_ALGN_EYE_IN_c;
input  RX_CLK_ALIGN_DONE_arst;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  debouncer_0_DB_OUT;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE;
output BIT_ALGN_ERR_0_c;
input  BIT_ALGN_OOR_c;
output BIT_ALGN_START_1_c;
output BIT_ALGN_DONE_c;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS;
input  PLL_LOCK_0;

    wire GND, VCC;
    
    
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_TRNG_Z1_1 
        u_CoreRxIODBitAlign (.BIT_ALGN_EYE_IN_c({BIT_ALGN_EYE_IN_c[2], 
        BIT_ALGN_EYE_IN_c[1], BIT_ALGN_EYE_IN_c[0]}), 
        .EYE_MONITOR_EARLY_net_0_0(EYE_MONITOR_EARLY_net_0_0), 
        .EYE_MONITOR_LATE_net_0_0(EYE_MONITOR_LATE_net_0_0), 
        .PLL_LOCK_0(PLL_LOCK_0), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS), .BIT_ALGN_DONE_c(
        BIT_ALGN_DONE_c), .BIT_ALGN_START_1_c(BIT_ALGN_START_1_c), 
        .BIT_ALGN_OOR_c(BIT_ALGN_OOR_c), .BIT_ALGN_ERR_0_c(
        BIT_ALGN_ERR_0_c), .CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module CORERXIODBITALIGN_C0_0(
       BIT_ALGN_EYE_IN_c,
       EYE_MONITOR_EARLY_net_0_0,
       EYE_MONITOR_LATE_net_0_0,
       PLL_LOCK_0,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS,
       BIT_ALGN_DONE_c,
       BIT_ALGN_START_1_c,
       BIT_ALGN_OOR_c,
       BIT_ALGN_ERR_0_c,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR,
       CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD,
       debouncer_0_DB_OUT,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst
    );
input  [2:0] BIT_ALGN_EYE_IN_c;
input  EYE_MONITOR_EARLY_net_0_0;
input  EYE_MONITOR_LATE_net_0_0;
input  PLL_LOCK_0;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS;
output BIT_ALGN_DONE_c;
output BIT_ALGN_START_1_c;
input  BIT_ALGN_OOR_c;
output BIT_ALGN_ERR_0_c;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR;
output CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD;
input  debouncer_0_DB_OUT;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  RX_CLK_ALIGN_DONE_arst;

    wire GND, VCC;
    
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
        CORERXIODBITALIGN_C0_CORERXIODBITALIGN_C0_0_CORERXIODBITALIGN_0s_0s_0s_26s_10s_10s_1 
        CORERXIODBITALIGN_C0_0 (.EYE_MONITOR_LATE_net_0_0(
        EYE_MONITOR_LATE_net_0_0), .EYE_MONITOR_EARLY_net_0_0(
        EYE_MONITOR_EARLY_net_0_0), .BIT_ALGN_EYE_IN_c({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE), .BIT_ALGN_ERR_0_c(
        BIT_ALGN_ERR_0_c), .BIT_ALGN_OOR_c(BIT_ALGN_OOR_c), 
        .BIT_ALGN_START_1_c(BIT_ALGN_START_1_c), .BIT_ALGN_DONE_c(
        BIT_ALGN_DONE_c), .CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS), .PLL_LOCK_0(
        PLL_LOCK_0));
    
endmodule


module PF_CCC_C0_PF_CCC_C0_0_PF_CCC(
       PF_OSC_C1_0_RCOSC_160MHZ_GL,
       PLL_LOCK_0,
       PF_CCC_C0_0_OUT0_FABCLK_0
    );
input  PF_OSC_C1_0_RCOSC_160MHZ_GL;
output PLL_LOCK_0;
output PF_CCC_C0_0_OUT0_FABCLK_0;

    wire [7:0] SSCG_WAVE_TABLE_ADDR_0;
    wire [32:0] DRI_RDATA_0;
    wire pll_inst_0_clkint_0, VCC, GND, DELAY_LINE_OUT_OF_RANGE_2, 
        OUT1, OUT2, OUT3, DRI_INTERRUPT_0;
    
    CLKINT clkint_0 (.A(pll_inst_0_clkint_0), .Y(
        PF_CCC_C0_0_OUT0_FABCLK_0));
    PLL #( .VCOFREQUENCY(5000), .DELAY_LINE_SIMULATION_MODE(""), .DATA_RATE(0.000000)
        , .FORMAL_NAME(""), .INTERFACE_NAME(""), .INTERFACE_LEVEL(32'b00000000000000000000000000000000)
        , .SOFTRESET(32'b00000000000000000000000000000000), .SOFT_POWERDOWN_N(32'b00000000000000000000000000000001)
        , .RFDIV_EN(32'b00000000000000000000000000000001), .OUT0_DIV_EN(32'b00000000000000000000000000000001)
        , .OUT1_DIV_EN(32'b00000000000000000000000000000000), .OUT2_DIV_EN(32'b00000000000000000000000000000000)
        , .OUT3_DIV_EN(32'b00000000000000000000000000000000), .SOFT_REF_CLK_SEL(32'b00000000000000000000000000000000)
        , .RESET_ON_LOCK(32'b00000000000000000000000000000001), .BYPASS_CLK_SEL(32'b00000000000000000000000000000000)
        , .BYPASS_GO_EN_N(32'b00000000000000000000000000000001), .BYPASS_PLL(32'b00000000000000000000000000000000)
        , .BYPASS_OUT_DIVIDER(32'b00000000000000000000000000000000), .FF_REQUIRES_LOCK(32'b00000000000000000000000000000000)
        , .FSE_N(32'b00000000000000000000000000000000), .FB_CLK_SEL_0(32'b00000000000000000000000000000000)
        , .FB_CLK_SEL_1(32'b00000000000000000000000000000000), .RFDIV(32'b00000000000000000000000000000100)
        , .FRAC_EN(32'b00000000000000000000000000000000), .FRAC_DAC_EN(32'b00000000000000000000000000000000)
        , .DIV0_RST_DELAY(32'b00000000000000000000000000000000), .DIV0_VAL(32'b00000000000000000000000000001010)
        , .DIV1_RST_DELAY(32'b00000000000000000000000000000000), .DIV1_VAL(32'b00000000000000000000000000000001)
        , .DIV2_RST_DELAY(32'b00000000000000000000000000000000), .DIV2_VAL(32'b00000000000000000000000000000001)
        , .DIV3_RST_DELAY(32'b00000000000000000000000000000000), .DIV3_VAL(32'b00000000000000000000000000000001)
        , .DIV3_CLK_SEL(32'b00000000000000000000000000000000), .BW_INT_CTRL(32'b00000000000000000000000000000000)
        , .BW_PROP_CTRL(32'b00000000000000000000000000000001), .IREF_EN(32'b00000000000000000000000000000001)
        , .IREF_TOGGLE(32'b00000000000000000000000000000000), .LOCK_CNT(32'b00000000000000000000000000001000)
        , .DESKEW_CAL_CNT(32'b00000000000000000000000000000110), .DESKEW_CAL_EN(32'b00000000000000000000000000000001)
        , .DESKEW_CAL_BYPASS(32'b00000000000000000000000000000000), .SYNC_REF_DIV_EN(32'b00000000000000000000000000000000)
        , .SYNC_REF_DIV_EN_2(32'b00000000000000000000000000000000), .OUT0_PHASE_SEL(32'b00000000000000000000000000000000)
        , .OUT1_PHASE_SEL(32'b00000000000000000000000000000000), .OUT2_PHASE_SEL(32'b00000000000000000000000000000000)
        , .OUT3_PHASE_SEL(32'b00000000000000000000000000000000), .SOFT_LOAD_PHASE_N(32'b00000000000000000000000000000001)
        , .SSM_DIV_VAL(32'b00000000000000000000000000000001), .FB_FRAC_VAL(32'b00000000000000000000000000000000)
        , .SSM_SPREAD_MODE(32'b00000000000000000000000000000000), .SSM_MODULATION(32'b00000000000000000000000000000101)
        , .FB_INT_VAL(32'b00000000000000000000000001111101), .SSM_EN_N(32'b00000000000000000000000000000001)
        , .SSM_EXT_WAVE_EN(32'b00000000000000000000000000000000), .SSM_EXT_WAVE_MAX_ADDR(32'b00000000000000000000000000000000)
        , .SSM_RANDOM_EN(32'b00000000000000000000000000000000), .SSM_RANDOM_PATTERN_SEL(32'b00000000000000000000000000000000)
        , .CDMUX0_SEL(32'b00000000000000000000000000000000), .CDMUX1_SEL(32'b00000000000000000000000000000001)
        , .CDMUX2_SEL(32'b00000000000000000000000000000000), .CDELAY0_SEL(32'b00000000000000000000000000000000)
        , .CDELAY0_EN(32'b00000000000000000000000000000000), .DRI_EN(32'b00000000000000000000000000000001)
         )  pll_inst_0 (.LOCK(PLL_LOCK_0), .SSCG_WAVE_TABLE_ADDR({
        SSCG_WAVE_TABLE_ADDR_0[7], SSCG_WAVE_TABLE_ADDR_0[6], 
        SSCG_WAVE_TABLE_ADDR_0[5], SSCG_WAVE_TABLE_ADDR_0[4], 
        SSCG_WAVE_TABLE_ADDR_0[3], SSCG_WAVE_TABLE_ADDR_0[2], 
        SSCG_WAVE_TABLE_ADDR_0[1], SSCG_WAVE_TABLE_ADDR_0[0]}), 
        .DELAY_LINE_OUT_OF_RANGE(DELAY_LINE_OUT_OF_RANGE_2), 
        .POWERDOWN_N(VCC), .OUT0_EN(VCC), .OUT1_EN(GND), .OUT2_EN(GND), 
        .OUT3_EN(GND), .REF_CLK_SEL(GND), .BYPASS_EN_N(VCC), 
        .LOAD_PHASE_N(VCC), .SSCG_WAVE_TABLE({GND, GND, GND, GND, GND, 
        GND, GND, GND}), .PHASE_DIRECTION(GND), .PHASE_ROTATE(GND), 
        .PHASE_OUT0_SEL(GND), .PHASE_OUT1_SEL(GND), .PHASE_OUT2_SEL(
        GND), .PHASE_OUT3_SEL(GND), .DELAY_LINE_MOVE(GND), 
        .DELAY_LINE_DIRECTION(GND), .DELAY_LINE_WIDE(GND), 
        .DELAY_LINE_LOAD(VCC), .REFCLK_SYNC_EN(GND), .REF_CLK_0(
        PF_OSC_C1_0_RCOSC_160MHZ_GL), .REF_CLK_1(GND), .FB_CLK(GND), 
        .OUT0(pll_inst_0_clkint_0), .OUT1(OUT1), .OUT2(OUT2), .OUT3(
        OUT3), .DRI_CLK(GND), .DRI_CTRL({GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .DRI_WDATA({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND}), .DRI_ARST_N(VCC), .DRI_RDATA({
        DRI_RDATA_0[32], DRI_RDATA_0[31], DRI_RDATA_0[30], 
        DRI_RDATA_0[29], DRI_RDATA_0[28], DRI_RDATA_0[27], 
        DRI_RDATA_0[26], DRI_RDATA_0[25], DRI_RDATA_0[24], 
        DRI_RDATA_0[23], DRI_RDATA_0[22], DRI_RDATA_0[21], 
        DRI_RDATA_0[20], DRI_RDATA_0[19], DRI_RDATA_0[18], 
        DRI_RDATA_0[17], DRI_RDATA_0[16], DRI_RDATA_0[15], 
        DRI_RDATA_0[14], DRI_RDATA_0[13], DRI_RDATA_0[12], 
        DRI_RDATA_0[11], DRI_RDATA_0[10], DRI_RDATA_0[9], 
        DRI_RDATA_0[8], DRI_RDATA_0[7], DRI_RDATA_0[6], DRI_RDATA_0[5], 
        DRI_RDATA_0[4], DRI_RDATA_0[3], DRI_RDATA_0[2], DRI_RDATA_0[1], 
        DRI_RDATA_0[0]}), .DRI_INTERRUPT(DRI_INTERRUPT_0));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule


module PF_CCC_C0(
       PF_CCC_C0_0_OUT0_FABCLK_0,
       PLL_LOCK_0,
       PF_OSC_C1_0_RCOSC_160MHZ_GL
    );
output PF_CCC_C0_0_OUT0_FABCLK_0;
output PLL_LOCK_0;
input  PF_OSC_C1_0_RCOSC_160MHZ_GL;

    wire GND, VCC;
    
    VCC VCC_Z (.Y(VCC));
    PF_CCC_C0_PF_CCC_C0_0_PF_CCC PF_CCC_C0_0 (
        .PF_OSC_C1_0_RCOSC_160MHZ_GL(PF_OSC_C1_0_RCOSC_160MHZ_GL), 
        .PLL_LOCK_0(PLL_LOCK_0), .PF_CCC_C0_0_OUT0_FABCLK_0(
        PF_CCC_C0_0_OUT0_FABCLK_0));
    GND GND_Z (.Y(GND));
    
endmodule


module ACT_UNIQUE_debouncer_1(
       SWITCH_c,
       PF_CCC_C0_0_OUT0_FABCLK_0,
       PLL_LOCK_0,
       DB_OUT_1z
    );
input  SWITCH_c;
input  PF_CCC_C0_0_OUT0_FABCLK_0;
input  PLL_LOCK_0;
output DB_OUT_1z;

    wire [3:0] q_reg_Z;
    wire [3:0] q_next_Z;
    wire VCC, DFF2_Z, GND, DFF1_Z, q_reset_Z, CO1;
    
    CFG3 #( .INIT(8'h20) )  \q_reg_RNI9STM[1]  (.A(q_reg_Z[0]), .B(
        q_reg_Z[3]), .C(q_reg_Z[1]), .Y(CO1));
    SLE DFF2 (.D(DFF1_Z), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), .EN(VCC), 
        .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(DFF2_Z));
    SLE DFF1 (.D(SWITCH_c), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), .EN(VCC), 
        .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(DFF1_Z));
    CFG3 #( .INIT(8'h12) )  \q_next[2]  (.A(q_reg_Z[2]), .B(q_reset_Z), 
        .C(CO1), .Y(q_next_Z[2]));
    GND GND_Z (.Y(GND));
    CFG2 #( .INIT(4'h6) )  q_reset (.A(DFF1_Z), .B(DFF2_Z), .Y(
        q_reset_Z));
    SLE \q_reg[2]  (.D(q_next_Z[2]), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), 
        .EN(VCC), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(q_reg_Z[2]));
    SLE \q_reg[0]  (.D(q_next_Z[0]), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), 
        .EN(VCC), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(q_reg_Z[0]));
    SLE \q_reg[1]  (.D(q_next_Z[1]), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), 
        .EN(VCC), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(q_reg_Z[1]));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'h006A) )  \q_next[3]  (.A(q_reg_Z[3]), .B(
        q_reg_Z[2]), .C(CO1), .D(q_reset_Z), .Y(q_next_Z[3]));
    CFG4 #( .INIT(16'h2130) )  \q_next[1]  (.A(q_reg_Z[3]), .B(
        q_reset_Z), .C(q_reg_Z[1]), .D(q_reg_Z[0]), .Y(q_next_Z[1]));
    SLE \q_reg[3]  (.D(q_next_Z[3]), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), 
        .EN(VCC), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(q_reg_Z[3]));
    SLE DB_OUT (.D(DFF2_Z), .CLK(PF_CCC_C0_0_OUT0_FABCLK_0), .EN(
        q_reg_Z[3]), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(DB_OUT_1z));
    CFG3 #( .INIT(8'h21) )  \q_next[0]  (.A(q_reg_Z[3]), .B(q_reset_Z), 
        .C(q_reg_Z[0]), .Y(q_next_Z[0]));
    
endmodule


module ACT_UNIQUE_prbscheck_parallel_fab_1(
       ACT_UNIQUE_rev_bits_0_out_data,
       prbs_chk_error_o_1_c,
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       RX_CLK_ALIGN_DONE_arst
    );
input  [7:0] ACT_UNIQUE_rev_bits_0_out_data;
output prbs_chk_error_o_1_c;
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  RX_CLK_ALIGN_DONE_arst;

    wire [6:0] s_in_old_Z;
    wire [7:0] s_error1_Z;
    wire [0:0] s_error1_2_Z;
    wire [1:1] s_error1_3_Z;
    wire [2:2] s_error1_4_Z;
    wire [3:3] s_error1_5_Z;
    wire [4:4] s_error1_6_Z;
    wire [5:5] s_error1_7_Z;
    wire [6:6] s_error1_8_Z;
    wire [7:7] s_error1_9_Z;
    wire VCC, GND, s_error0_Z, un1_s_error0_i, s_prbs_chk_error_Z, 
        un1_s_error0_4_Z, s_prbs_chk_error_5_Z, s_prbs_chk_error_4_Z;
    
    CFG3 #( .INIT(8'h96) )  \s_error1_8[6]  (.A(s_in_old_Z[4]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[6]), .C(s_in_old_Z[5]), .Y(
        s_error1_8_Z[6]));
    GND GND_Z (.Y(GND));
    SLE \s_in_old[0]  (.D(ACT_UNIQUE_rev_bits_0_out_data[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[0]));
    CFG4 #( .INIT(16'hFFFE) )  un1_s_error0_4 (.A(
        ACT_UNIQUE_rev_bits_0_out_data[3]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[1]), .C(
        ACT_UNIQUE_rev_bits_0_out_data[2]), .D(
        ACT_UNIQUE_rev_bits_0_out_data[6]), .Y(un1_s_error0_4_Z));
    SLE \s_in_old[6]  (.D(ACT_UNIQUE_rev_bits_0_out_data[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[6]));
    SLE \s_in_old[3]  (.D(ACT_UNIQUE_rev_bits_0_out_data[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[3]));
    SLE \s_error1[7]  (.D(s_error1_9_Z[7]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[7]));
    VCC VCC_Z (.Y(VCC));
    SLE \s_error1[6]  (.D(s_error1_8_Z[6]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[6]));
    SLE prbs_chk_error_o (.D(s_prbs_chk_error_Z), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(prbs_chk_error_o_1_c));
    SLE \s_error1[0]  (.D(s_error1_2_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[0]));
    CFG3 #( .INIT(8'h96) )  \s_error1_6[4]  (.A(s_in_old_Z[2]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[4]), .C(s_in_old_Z[3]), .Y(
        s_error1_6_Z[4]));
    CFG3 #( .INIT(8'h96) )  \s_error1_5[3]  (.A(s_in_old_Z[1]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[3]), .C(s_in_old_Z[2]), .Y(
        s_error1_5_Z[3]));
    SLE \s_error1[1]  (.D(s_error1_3_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[1]));
    CFG4 #( .INIT(16'hFFFE) )  s_prbs_chk_error (.A(s_error1_Z[4]), .B(
        s_error1_Z[5]), .C(s_prbs_chk_error_5_Z), .D(
        s_prbs_chk_error_4_Z), .Y(s_prbs_chk_error_Z));
    SLE \s_in_old[1]  (.D(ACT_UNIQUE_rev_bits_0_out_data[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[1]));
    CFG4 #( .INIT(16'hFFFE) )  s_prbs_chk_error_5 (.A(s_error1_Z[3]), 
        .B(s_error1_Z[2]), .C(s_error1_Z[1]), .D(s_error1_Z[0]), .Y(
        s_prbs_chk_error_5_Z));
    SLE \s_error1[3]  (.D(s_error1_5_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[3]));
    SLE \s_in_old[4]  (.D(ACT_UNIQUE_rev_bits_0_out_data[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[4]));
    CFG3 #( .INIT(8'h96) )  \s_error1_9[7]  (.A(s_in_old_Z[5]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[7]), .C(s_in_old_Z[6]), .Y(
        s_error1_9_Z[7]));
    CFG3 #( .INIT(8'h96) )  \s_error1_2[0]  (.A(
        ACT_UNIQUE_rev_bits_0_out_data[6]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[7]), .C(
        ACT_UNIQUE_rev_bits_0_out_data[0]), .Y(s_error1_2_Z[0]));
    SLE \s_in_old[5]  (.D(ACT_UNIQUE_rev_bits_0_out_data[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[5]));
    SLE \s_error1[2]  (.D(s_error1_4_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[2]));
    CFG4 #( .INIT(16'h0001) )  s_error0_RNO (.A(
        ACT_UNIQUE_rev_bits_0_out_data[5]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[0]), .C(
        ACT_UNIQUE_rev_bits_0_out_data[4]), .D(un1_s_error0_4_Z), .Y(
        un1_s_error0_i));
    SLE s_error0 (.D(un1_s_error0_i), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error0_Z));
    SLE \s_in_old[2]  (.D(ACT_UNIQUE_rev_bits_0_out_data[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_in_old_Z[2]));
    CFG3 #( .INIT(8'h96) )  \s_error1_3[1]  (.A(
        ACT_UNIQUE_rev_bits_0_out_data[1]), .B(s_in_old_Z[0]), .C(
        ACT_UNIQUE_rev_bits_0_out_data[7]), .Y(s_error1_3_Z[1]));
    CFG3 #( .INIT(8'h96) )  \s_error1_4[2]  (.A(s_in_old_Z[0]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[2]), .C(s_in_old_Z[1]), .Y(
        s_error1_4_Z[2]));
    CFG3 #( .INIT(8'h96) )  \s_error1_7[5]  (.A(s_in_old_Z[3]), .B(
        ACT_UNIQUE_rev_bits_0_out_data[5]), .C(s_in_old_Z[4]), .Y(
        s_error1_7_Z[5]));
    SLE \s_error1[5]  (.D(s_error1_7_Z[5]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[5]));
    CFG3 #( .INIT(8'hFE) )  s_prbs_chk_error_4 (.A(s_error1_Z[7]), .B(
        s_error1_Z[6]), .C(s_error0_Z), .Y(s_prbs_chk_error_4_Z));
    SLE \s_error1[4]  (.D(s_error1_6_Z[4]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(
        RX_CLK_ALIGN_DONE_arst), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(s_error1_Z[4]));
    
endmodule


module ACT_UNIQUE_debouncer_0(
       PF_IOD_GENERIC_RX_C1_0_RX_CLK_G,
       PLL_LOCK_0,
       debouncer_0_DB_OUT,
       RESTARTN_c
    );
input  PF_IOD_GENERIC_RX_C1_0_RX_CLK_G;
input  PLL_LOCK_0;
output debouncer_0_DB_OUT;
input  RESTARTN_c;

    wire [3:0] q_reg_Z;
    wire [3:0] q_next_Z;
    wire RESTARTN_c_i, VCC, DFF2_Z, GND, DFF1_Z, q_reset_0, CO1;
    
    SLE DFF2 (.D(DFF1_Z), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        VCC), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(DFF2_Z));
    SLE DFF1 (.D(RESTARTN_c_i), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), 
        .EN(VCC), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(DFF1_Z));
    CFG3 #( .INIT(8'h12) )  \q_next[2]  (.A(q_reg_Z[2]), .B(q_reset_0), 
        .C(CO1), .Y(q_next_Z[2]));
    GND GND_Z (.Y(GND));
    CFG2 #( .INIT(4'h6) )  q_reset (.A(DFF1_Z), .B(DFF2_Z), .Y(
        q_reset_0));
    CFG3 #( .INIT(8'h20) )  \q_reg_RNI26281[1]  (.A(q_reg_Z[0]), .B(
        q_reg_Z[3]), .C(q_reg_Z[1]), .Y(CO1));
    SLE \q_reg[2]  (.D(q_next_Z[2]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(PLL_LOCK_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(q_reg_Z[2]));
    SLE \q_reg[0]  (.D(q_next_Z[0]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(PLL_LOCK_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(q_reg_Z[0]));
    SLE \q_reg[1]  (.D(q_next_Z[1]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(PLL_LOCK_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(q_reg_Z[1]));
    VCC VCC_Z (.Y(VCC));
    CFG4 #( .INIT(16'h006A) )  \q_next[3]  (.A(q_reg_Z[3]), .B(
        q_reg_Z[2]), .C(CO1), .D(q_reset_0), .Y(q_next_Z[3]));
    CFG1 #( .INIT(2'h1) )  DFF1_RNO (.A(RESTARTN_c), .Y(RESTARTN_c_i));
    CFG4 #( .INIT(16'h2130) )  \q_next[1]  (.A(q_reg_Z[3]), .B(
        q_reset_0), .C(q_reg_Z[1]), .D(q_reg_Z[0]), .Y(q_next_Z[1]));
    SLE \q_reg[3]  (.D(q_next_Z[3]), .CLK(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(VCC), .ALn(PLL_LOCK_0), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(q_reg_Z[3]));
    SLE DB_OUT (.D(DFF2_Z), .CLK(PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .EN(
        q_reg_Z[3]), .ALn(PLL_LOCK_0), .ADn(VCC), .SLn(VCC), .SD(GND), 
        .LAT(GND), .Q(debouncer_0_DB_OUT));
    CFG3 #( .INIT(8'h21) )  \q_next[0]  (.A(q_reg_Z[3]), .B(q_reset_0), 
        .C(q_reg_Z[0]), .Y(q_next_Z[0]));
    
endmodule


module IOG_IOD_DDRX4_COMP(
       BIT_ALGN_EYE_IN,
       RESTARTN,
       RXD,
       RXD_N,
       RX_CLK_N,
       RX_CLK_P,
       SWITCH,
       Algn_Done,
       Algn_Err,
       BIT_ALGN_DONE,
       BIT_ALGN_DONE_0,
       BIT_ALGN_ERR,
       BIT_ALGN_ERR_0,
       BIT_ALGN_OOR,
       BIT_ALGN_OOR_0,
       BIT_ALGN_START,
       BIT_ALGN_START_0,
       BIT_ALGN_START_1,
       CLK_TRAIN_ERROR,
       PLL_LOCK,
       PLL_LOCK_0,
       PRBS_ERR,
       PRBS_ERR_0,
       TXD,
       TXD_N,
       TX_CLK,
       TX_CLK_N,
       Y,
       prbs_chk_error_o_1
    );
input  [2:0] BIT_ALGN_EYE_IN;
input  RESTARTN;
input  [1:0] RXD;
input  [1:0] RXD_N;
input  RX_CLK_N;
input  RX_CLK_P;
input  SWITCH;
output Algn_Done;
output Algn_Err;
output BIT_ALGN_DONE;
output BIT_ALGN_DONE_0;
output BIT_ALGN_ERR;
output BIT_ALGN_ERR_0;
output BIT_ALGN_OOR;
output BIT_ALGN_OOR_0;
output BIT_ALGN_START;
output BIT_ALGN_START_0;
output BIT_ALGN_START_1;
output CLK_TRAIN_ERROR;
output PLL_LOCK;
output PLL_LOCK_0;
output PRBS_ERR;
output PRBS_ERR_0;
output [1:0] TXD;
output [1:0] TXD_N;
output TX_CLK;
output TX_CLK_N;
output Y;
output prbs_chk_error_o_1;

    wire [7:0] ACT_UNIQUE_rev_bits_0_out_data;
    wire [1:0] EYE_MONITOR_EARLY_net_0;
    wire [1:0] EYE_MONITOR_LATE_net_0;
    wire [7:0] rev_bits_0_out_data_4;
    wire [7:0] prbsgen_parallel_fab_0_prbs_out_msb_o_0;
    wire [3:0] PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX;
    wire [2:0] 
        \CORERXIODBITALIGN_C0_1.CORERXIODBITALIGN_C0_0.rx_BIT_ALGN_EYE_OUT ;
    wire [2:0] 
        \CORERXIODBITALIGN_C0_0.CORERXIODBITALIGN_C0_0.rx_BIT_ALGN_EYE_OUT ;
    wire [7:7] 
        \PF_IOD_TX_CCC_C0_0.COREBCLKSCLKALIGN_0.PF_IOD_TX_CCC_C0_TR_0.genblk1.U_PLL_BCLKSCLKALIGN.current_state ;
    wire [2:0] BIT_ALGN_EYE_IN_c;
    wire [7:0] \PF_IOD_GENERIC_RX_C1_0.un1_COREBCLKSCLKALIGN_0 ;
    wire [7:0] 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.ICB_CLK_ALGN_TAPDLY ;
    wire [7:0] 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.PF_IOD_GENERIC_RX_C1_TR_0.ICB_CLK_ALGN_TAPDLY ;
    wire PF_CCC_C0_0_OUT0_FABCLK_0, PF_IOD_GENERIC_RX_C1_0_RX_CLK_G, 
        debouncer_0_DB_OUT, CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS, 
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR, 
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD, 
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE, 
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS, 
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR, 
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD, 
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE, 
        PF_OSC_C1_0_RCOSC_160MHZ_GL, 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0, 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90, 
        PF_IOD_TX_CCC_C0_0_TX_CLK_G, VCC, GND, RX_CLK_ALIGN_DONE_arst, 
        \CORERXIODBITALIGN_C0_1.CORERXIODBITALIGN_C0_0.popfeedthru_unused , 
        \CORERXIODBITALIGN_C0_0.CORERXIODBITALIGN_C0_0.popfeedthru_unused , 
        \PF_CCC_C0_0.PF_CCC_C0_0.PLL_LOCK_0 , 
        \PF_IOD_TX_CCC_C0_0.PF_CCC_0.PLL_LOCK_0 , 
        \ACT_UNIQUE_debouncer_0.DB_OUT , N_81, RESTARTN_c, SWITCH_c, 
        BIT_ALGN_DONE_c, BIT_ALGN_DONE_0_c, BIT_ALGN_ERR_c, 
        BIT_ALGN_ERR_0_c, BIT_ALGN_OOR_c, BIT_ALGN_OOR_0_c, 
        BIT_ALGN_START_0_c, BIT_ALGN_START_1_c, CLK_TRAIN_ERROR_c, 
        PRBS_ERR_0_c, Y_c, prbs_chk_error_o_1_c, PLL_LOCK_c_i, 
        \PF_IOD_GENERIC_RX_C1_0.N_1 , \PF_IOD_GENERIC_RX_C1_0.N_2 , 
        \PF_IOD_GENERIC_RX_C1_0.N_3 , \PF_IOD_GENERIC_RX_C1_0.N_4 , 
        \PF_IOD_GENERIC_RX_C1_0.N_5 , \PF_IOD_GENERIC_RX_C1_0.N_6 , 
        \PF_IOD_GENERIC_RX_C1_0.N_7 , \PF_IOD_GENERIC_RX_C1_0.N_8 , 
        \PF_IOD_GENERIC_RX_C1_0.N_9 , \PF_IOD_GENERIC_RX_C1_0.N_10 , 
        \PF_IOD_GENERIC_RX_C1_0.N_11 , \PF_IOD_GENERIC_RX_C1_0.N_12 , 
        \PF_IOD_GENERIC_RX_C1_0.N_13 , \PF_IOD_GENERIC_RX_C1_0.N_14 , 
        \PF_IOD_GENERIC_RX_C1_0.N_16 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_1 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_2 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_3 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_4 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_5 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_6 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_7 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_8 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_9 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_10 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_11 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_12 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_13 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_14 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.N_33 , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.PF_IOD_GENERIC_RX_C1_TR_0.genblk1.un1_U_ICB_BCLKSCLKALIGN , 
        \PF_IOD_GENERIC_RX_C1_0.COREBCLKSCLKALIGN_0.PF_IOD_GENERIC_RX_C1_TR_0.N_1 ;
    
    INBUF SWITCH_ibuf (.PAD(SWITCH), .Y(SWITCH_c));
    ACT_UNIQUE_prbsgen_parallel_fab prbsgen_parallel_fab_0 (
        .prbsgen_parallel_fab_0_prbs_out_msb_o_0({
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[0]}), .current_state_0(
        \PF_IOD_TX_CCC_C0_0.COREBCLKSCLKALIGN_0.PF_IOD_TX_CCC_C0_TR_0.genblk1.U_PLL_BCLKSCLKALIGN.current_state [7])
        , .PF_IOD_TX_CCC_C0_0_TX_CLK_G(PF_IOD_TX_CCC_C0_0_TX_CLK_G));
    INBUF \BIT_ALGN_EYE_IN_ibuf[0]  (.PAD(BIT_ALGN_EYE_IN[0]), .Y(
        BIT_ALGN_EYE_IN_c[0]));
    PF_IOD_TX_CCC_C0 PF_IOD_TX_CCC_C0_0 (
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX({
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]}), 
        .current_state_0(
        \PF_IOD_TX_CCC_C0_0.COREBCLKSCLKALIGN_0.PF_IOD_TX_CCC_C0_TR_0.genblk1.U_PLL_BCLKSCLKALIGN.current_state [7])
        , .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0), .PLL_LOCK_c_i(
        PLL_LOCK_c_i), .PF_CCC_C0_0_OUT0_FABCLK_0(
        PF_CCC_C0_0_OUT0_FABCLK_0), .DB_OUT(
        \ACT_UNIQUE_debouncer_0.DB_OUT ), .PF_IOD_TX_CCC_C0_0_TX_CLK_G(
        PF_IOD_TX_CCC_C0_0_TX_CLK_G), .N_81(N_81), .PLL_LOCK_0(
        \PF_IOD_TX_CCC_C0_0.PF_CCC_0.PLL_LOCK_0 ));
    OUTBUF BIT_ALGN_START_1_obuf (.D(BIT_ALGN_START_1_c), .PAD(
        BIT_ALGN_START_1));
    OUTBUF Algn_Err_obuf (.D(BIT_ALGN_ERR_c), .PAD(Algn_Err));
    BUFF BUFF_0 (.A(RESTARTN_c), .Y(Y_c));
    ACT_UNIQUE_prbscheck_parallel_fab 
        ACT_UNIQUE_prbscheck_parallel_fab_0 (.rev_bits_0_out_data_4({
        rev_bits_0_out_data_4[7], rev_bits_0_out_data_4[6], 
        rev_bits_0_out_data_4[5], rev_bits_0_out_data_4[4], 
        rev_bits_0_out_data_4[3], rev_bits_0_out_data_4[2], 
        rev_bits_0_out_data_4[1], rev_bits_0_out_data_4[0]}), 
        .PRBS_ERR_0_c(PRBS_ERR_0_c), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst));
    INBUF RESTARTN_ibuf (.PAD(RESTARTN), .Y(RESTARTN_c));
    OUTBUF PLL_LOCK_obuf (.D(\PF_IOD_TX_CCC_C0_0.PF_CCC_0.PLL_LOCK_0 ), 
        .PAD(PLL_LOCK));
    INBUF \BIT_ALGN_EYE_IN_ibuf[1]  (.PAD(BIT_ALGN_EYE_IN[1]), .Y(
        BIT_ALGN_EYE_IN_c[1]));
    PF_IOD_GENERIC_RX_C1 PF_IOD_GENERIC_RX_C1_0 (.BIT_ALGN_EYE_IN_c({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .RXD_N({RXD_N[1], RXD_N[0]}), .RXD({
        RXD[1], RXD[0]}), .rev_bits_0_out_data_4({
        rev_bits_0_out_data_4[7], rev_bits_0_out_data_4[6], 
        rev_bits_0_out_data_4[5], rev_bits_0_out_data_4[4], 
        rev_bits_0_out_data_4[3], rev_bits_0_out_data_4[2], 
        rev_bits_0_out_data_4[1], rev_bits_0_out_data_4[0]}), 
        .EYE_MONITOR_EARLY_net_0({EYE_MONITOR_EARLY_net_0[1], 
        EYE_MONITOR_EARLY_net_0[0]}), .EYE_MONITOR_LATE_net_0({
        EYE_MONITOR_LATE_net_0[1], EYE_MONITOR_LATE_net_0[0]}), 
        .ACT_UNIQUE_rev_bits_0_out_data({
        ACT_UNIQUE_rev_bits_0_out_data[7], 
        ACT_UNIQUE_rev_bits_0_out_data[6], 
        ACT_UNIQUE_rev_bits_0_out_data[5], 
        ACT_UNIQUE_rev_bits_0_out_data[4], 
        ACT_UNIQUE_rev_bits_0_out_data[3], 
        ACT_UNIQUE_rev_bits_0_out_data[2], 
        ACT_UNIQUE_rev_bits_0_out_data[1], 
        ACT_UNIQUE_rev_bits_0_out_data[0]}), .current_state_0(
        \PF_IOD_TX_CCC_C0_0.COREBCLKSCLKALIGN_0.PF_IOD_TX_CCC_C0_TR_0.genblk1.U_PLL_BCLKSCLKALIGN.current_state [7])
        , .CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD), .BIT_ALGN_OOR_0_c(
        BIT_ALGN_OOR_0_c), .CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD), .BIT_ALGN_OOR_c(
        BIT_ALGN_OOR_c), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst), .CLK_TRAIN_ERROR_c(CLK_TRAIN_ERROR_c), 
        .RX_CLK_P(RX_CLK_P), .RX_CLK_N(RX_CLK_N), 
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G));
    CORERXIODBITALIGN_C0_1 CORERXIODBITALIGN_C0_0 (.BIT_ALGN_EYE_IN_c({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .EYE_MONITOR_EARLY_net_0_0(
        EYE_MONITOR_EARLY_net_0[0]), .EYE_MONITOR_LATE_net_0_0(
        EYE_MONITOR_LATE_net_0[0]), .PLL_LOCK_0(
        \PF_IOD_TX_CCC_C0_0.PF_CCC_0.PLL_LOCK_0 ), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_CLR_FLGS), .BIT_ALGN_DONE_0_c(
        BIT_ALGN_DONE_0_c), .BIT_ALGN_START_0_c(BIT_ALGN_START_0_c), 
        .BIT_ALGN_OOR_0_c(BIT_ALGN_OOR_0_c), .BIT_ALGN_ERR_c(
        BIT_ALGN_ERR_c), .CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_0_BIT_ALGN_LOAD), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst));
    OUTBUF PLL_LOCK_0_obuf (.D(\PF_CCC_C0_0.PF_CCC_C0_0.PLL_LOCK_0 ), 
        .PAD(PLL_LOCK_0));
    OUTBUF BIT_ALGN_DONE_obuf (.D(BIT_ALGN_DONE_c), .PAD(BIT_ALGN_DONE)
        );
    OUTBUF BIT_ALGN_START_0_obuf (.D(BIT_ALGN_START_0_c), .PAD(
        BIT_ALGN_START_0));
    OUTBUF Y_obuf (.D(Y_c), .PAD(Y));
    OUTBUF prbs_chk_error_o_1_obuf (.D(prbs_chk_error_o_1_c), .PAD(
        prbs_chk_error_o_1));
    INBUF \BIT_ALGN_EYE_IN_ibuf[2]  (.PAD(BIT_ALGN_EYE_IN[2]), .Y(
        BIT_ALGN_EYE_IN_c[2]));
    PF_OSC_C1 PF_OSC_C1_0 (.PF_OSC_C1_0_RCOSC_160MHZ_GL(
        PF_OSC_C1_0_RCOSC_160MHZ_GL));
    PF_IOD_GENERIC_TX_C0 PF_IOD_GENERIC_TX_C0_0 (
        .prbsgen_parallel_fab_0_prbs_out_msb_o_0({
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[7], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[6], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[5], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[4], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[3], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[2], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[1], 
        prbsgen_parallel_fab_0_prbs_out_msb_o_0[0]}), .TXD_N({TXD_N[1], 
        TXD_N[0]}), .TXD({TXD[1], TXD[0]}), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX({
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[3], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[2], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[1], 
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_CLK_ALIGN_IOD_RX[0]}), 
        .TX_CLK_N(TX_CLK_N), .TX_CLK(TX_CLK), 
        .PF_IOD_TX_CCC_C0_0_TX_CLK_G(PF_IOD_TX_CCC_C0_0_TX_CLK_G), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_90), 
        .PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0(
        PF_IOD_TX_CCC_C0_0_IOD_TX_CLKS_HS_IO_CLK_0), .PLL_LOCK_c_i(
        PLL_LOCK_c_i), .N_81(N_81));
    OUTBUF PRBS_ERR_obuf (.D(PRBS_ERR_0_c), .PAD(PRBS_ERR));
    OUTBUF BIT_ALGN_OOR_0_obuf (.D(BIT_ALGN_OOR_0_c), .PAD(
        BIT_ALGN_OOR_0));
    GND GND_Z (.Y(GND));
    OUTBUF BIT_ALGN_ERR_obuf (.D(BIT_ALGN_ERR_c), .PAD(BIT_ALGN_ERR));
    VCC VCC_Z (.Y(VCC));
    CORERXIODBITALIGN_C0_0 CORERXIODBITALIGN_C0_1 (.BIT_ALGN_EYE_IN_c({
        BIT_ALGN_EYE_IN_c[2], BIT_ALGN_EYE_IN_c[1], 
        BIT_ALGN_EYE_IN_c[0]}), .EYE_MONITOR_EARLY_net_0_0(
        EYE_MONITOR_EARLY_net_0[1]), .EYE_MONITOR_LATE_net_0_0(
        EYE_MONITOR_LATE_net_0[1]), .PLL_LOCK_0(
        \PF_IOD_TX_CCC_C0_0.PF_CCC_0.PLL_LOCK_0 ), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_CLR_FLGS), .BIT_ALGN_DONE_c(
        BIT_ALGN_DONE_c), .BIT_ALGN_START_1_c(BIT_ALGN_START_1_c), 
        .BIT_ALGN_OOR_c(BIT_ALGN_OOR_c), .BIT_ALGN_ERR_0_c(
        BIT_ALGN_ERR_0_c), .CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_MOVE), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_DIR), 
        .CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD(
        CORERXIODBITALIGN_C0_1_BIT_ALGN_LOAD), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst));
    OUTBUF PRBS_ERR_0_obuf (.D(PRBS_ERR_0_c), .PAD(PRBS_ERR_0));
    PF_CCC_C0 PF_CCC_C0_0 (.PF_CCC_C0_0_OUT0_FABCLK_0(
        PF_CCC_C0_0_OUT0_FABCLK_0), .PLL_LOCK_0(
        \PF_CCC_C0_0.PF_CCC_C0_0.PLL_LOCK_0 ), 
        .PF_OSC_C1_0_RCOSC_160MHZ_GL(PF_OSC_C1_0_RCOSC_160MHZ_GL));
    OUTBUF BIT_ALGN_DONE_0_obuf (.D(BIT_ALGN_DONE_0_c), .PAD(
        BIT_ALGN_DONE_0));
    ACT_UNIQUE_debouncer_1 ACT_UNIQUE_debouncer_0 (.SWITCH_c(SWITCH_c), 
        .PF_CCC_C0_0_OUT0_FABCLK_0(PF_CCC_C0_0_OUT0_FABCLK_0), 
        .PLL_LOCK_0(\PF_CCC_C0_0.PF_CCC_C0_0.PLL_LOCK_0 ), .DB_OUT_1z(
        \ACT_UNIQUE_debouncer_0.DB_OUT ));
    OUTBUF CLK_TRAIN_ERROR_obuf (.D(CLK_TRAIN_ERROR_c), .PAD(
        CLK_TRAIN_ERROR));
    OUTBUF Algn_Done_obuf (.D(BIT_ALGN_DONE_0_c), .PAD(Algn_Done));
    OUTBUF BIT_ALGN_START_obuf (.D(BIT_ALGN_START_0_c), .PAD(
        BIT_ALGN_START));
    ACT_UNIQUE_prbscheck_parallel_fab_1 
        ACT_UNIQUE_prbscheck_parallel_fab_1 (
        .ACT_UNIQUE_rev_bits_0_out_data({
        ACT_UNIQUE_rev_bits_0_out_data[7], 
        ACT_UNIQUE_rev_bits_0_out_data[6], 
        ACT_UNIQUE_rev_bits_0_out_data[5], 
        ACT_UNIQUE_rev_bits_0_out_data[4], 
        ACT_UNIQUE_rev_bits_0_out_data[3], 
        ACT_UNIQUE_rev_bits_0_out_data[2], 
        ACT_UNIQUE_rev_bits_0_out_data[1], 
        ACT_UNIQUE_rev_bits_0_out_data[0]}), .prbs_chk_error_o_1_c(
        prbs_chk_error_o_1_c), .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .RX_CLK_ALIGN_DONE_arst(
        RX_CLK_ALIGN_DONE_arst));
    OUTBUF BIT_ALGN_ERR_0_obuf (.D(BIT_ALGN_ERR_0_c), .PAD(
        BIT_ALGN_ERR_0));
    ACT_UNIQUE_debouncer_0 debouncer_0 (
        .PF_IOD_GENERIC_RX_C1_0_RX_CLK_G(
        PF_IOD_GENERIC_RX_C1_0_RX_CLK_G), .PLL_LOCK_0(
        \PF_IOD_TX_CCC_C0_0.PF_CCC_0.PLL_LOCK_0 ), .debouncer_0_DB_OUT(
        debouncer_0_DB_OUT), .RESTARTN_c(RESTARTN_c));
    OUTBUF BIT_ALGN_OOR_obuf (.D(BIT_ALGN_OOR_c), .PAD(BIT_ALGN_OOR));
    
endmodule
