// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAI110I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAlOlOI
,
CAXI4DMAIOlOI
,
CAXI4DMAllI0I
,
CAXI4DMAl0IlI
,
CAXI4DMAI0I0I
)
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAlOlOI
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAIOlOI
;
input
CAXI4DMAllI0I
;
output
CAXI4DMAl0IlI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0I0I
;
reg
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAl101I
;
wire
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOO11I
;
wire
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAIO11I
;
integer
CAXI4DMAlO11I
;
wire
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAIlO0I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl101I
<=
{
NUM_INT_BDS
{
1
'b
0
}
}
;
end
else
begin
for
(
CAXI4DMAlO11I
=
0
;
CAXI4DMAlO11I
<
NUM_INT_BDS
;
CAXI4DMAlO11I
=
CAXI4DMAlO11I
+
1
)
begin
if
(
CAXI4DMAOO11I
[
CAXI4DMAlO11I
]
)
begin
CAXI4DMAl101I
[
CAXI4DMAlO11I
]
<=
1
'b
1
;
end
else
if
(
CAXI4DMAIO11I
[
CAXI4DMAlO11I
]
)
begin
CAXI4DMAl101I
[
CAXI4DMAlO11I
]
<=
1
'b
0
;
end
end
end
end
CAXI4DMAOI11I
#
(
.CAXI4DMAIl1lI
(
NUM_INT_BDS
)
)
CAXI4DMAII11I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO01lI
(
CAXI4DMAl101I
)
,
.CAXI4DMAlI11I
(
CAXI4DMAllI0I
)
,
.CAXI4DMAOl11I
(
CAXI4DMAIO11I
)
,
.CAXI4DMAIlO0I
(
CAXI4DMAIlO0I
)
)
;
assign
CAXI4DMAOO11I
=
CAXI4DMAlOlOI
|
CAXI4DMAIOlOI
;
assign
CAXI4DMAI0I0I
=
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000000000010
)
?
'd
1
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000000000100
)
?
'd
2
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000000001000
)
?
'd
3
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000000010000
)
?
'd
4
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000000100000
)
?
'd
5
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000001000000
)
?
'd
6
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000010000000
)
?
'd
7
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000000100000000
)
?
'd
8
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000001000000000
)
?
'd
9
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000010000000000
)
?
'd
10
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000000100000000000
)
?
'd
11
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000001000000000000
)
?
'd
12
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000010000000000000
)
?
'd
13
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000000100000000000000
)
?
'd
14
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000001000000000000000
)
?
'd
15
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000010000000000000000
)
?
'd
16
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000000100000000000000000
)
?
'd
17
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000001000000000000000000
)
?
'd
18
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000010000000000000000000
)
?
'd
19
:
(
CAXI4DMAIlO0I
==
32
'b
00000000000100000000000000000000
)
?
'd
20
:
(
CAXI4DMAIlO0I
==
32
'b
00000000001000000000000000000000
)
?
'd
21
:
(
CAXI4DMAIlO0I
==
32
'b
00000000010000000000000000000000
)
?
'd
22
:
(
CAXI4DMAIlO0I
==
32
'b
00000000100000000000000000000000
)
?
'd
23
:
(
CAXI4DMAIlO0I
==
32
'b
00000001000000000000000000000000
)
?
'd
24
:
(
CAXI4DMAIlO0I
==
32
'b
00000010000000000000000000000000
)
?
'd
25
:
(
CAXI4DMAIlO0I
==
32
'b
00000100000000000000000000000000
)
?
'd
26
:
(
CAXI4DMAIlO0I
==
32
'b
00001000000000000000000000000000
)
?
'd
27
:
(
CAXI4DMAIlO0I
==
32
'b
00010000000000000000000000000000
)
?
'd
28
:
(
CAXI4DMAIlO0I
==
32
'b
00100000000000000000000000000000
)
?
'd
29
:
(
CAXI4DMAIlO0I
==
32
'b
01000000000000000000000000000000
)
?
'd
30
:
(
CAXI4DMAIlO0I
==
32
'b
10000000000000000000000000000000
)
?
'd
31
:
'd
0
;
assign
CAXI4DMAl0IlI
=
(
|
CAXI4DMAIlO0I
)
;
endmodule
