//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Oct  7 17:23:30 2020
// Version: v12.4 12.900.0.16
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// Top
module Top(
    // Inputs
    CLK_0,
    D,
    // Outputs
    Q
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  CLK_0;
input  D;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Q;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   CLK_0;
wire   D;
wire   DFN1_0_Q;
wire   DFN1_1_Q;
wire   Q_net_0;
wire   Q_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Q_net_1 = Q_net_0;
assign Q       = Q_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------DFN1
DFN1 DFN1_0(
        // Inputs
        .D   ( D ),
        .CLK ( CLK_0 ),
        // Outputs
        .Q   ( DFN1_0_Q ) 
        );

//--------DFN1
DFN1 DFN1_1(
        // Inputs
        .D   ( DFN1_0_Q ),
        .CLK ( CLK_0 ),
        // Outputs
        .Q   ( DFN1_1_Q ) 
        );

//--------DFN1
DFN1 DFN1_2(
        // Inputs
        .D   ( DFN1_1_Q ),
        .CLK ( CLK_0 ),
        // Outputs
        .Q   ( Q_net_0 ) 
        );


endmodule
