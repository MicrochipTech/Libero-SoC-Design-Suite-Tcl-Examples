// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAIIO0I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAO01lI
,
CAXI4DMAOlO0I
,
CAXI4DMAIlO0I
)
;
parameter
CAXI4DMAIl1lI
=
4
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAO01lI
;
input
CAXI4DMAOlO0I
;
output
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAIlO0I
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAO1O1l
;
reg
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAI1O1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAl1O1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAOOI1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAIOI1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAlOI1l
;
assign
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
1
:
0
]
&
CAXI4DMAI1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
assign
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
1
:
1
]
=
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
2
:
0
]
|
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
2
:
0
]
;
assign
CAXI4DMAl1O1l
[
0
]
=
1
'b
0
;
assign
CAXI4DMAOOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
&
~
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
assign
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
1
:
1
]
=
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
2
:
0
]
|
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
2
:
0
]
;
assign
CAXI4DMAIOI1l
[
0
]
=
1
'b
0
;
assign
CAXI4DMAlOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
1
:
0
]
&
~
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
assign
CAXI4DMAIlO0I
[
CAXI4DMAIl1lI
-
1
:
0
]
=
(
|
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
)
?
CAXI4DMAOOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
:
CAXI4DMAlOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1O1l
<=
{
CAXI4DMAIl1lI
{
1
'b
1
}
}
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
if
(
|
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
)
begin
CAXI4DMAI1O1l
<=
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
end
else
begin
CAXI4DMAI1O1l
<=
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
end
end
end
endmodule
