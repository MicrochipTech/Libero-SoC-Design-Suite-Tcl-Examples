// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAl1IOI
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAIOlOI
,
CAXI4DMAlOlOI
,
CAXI4DMAI1l
,
CAXI4DMAl1l
,
CAXI4DMAOO0
,
CAXI4DMAIO0
,
CAXI4DMAlO0
,
CAXI4DMAOI0
,
CAXI4DMAII0
,
CAXI4DMAlI0
,
CAXI4DMAOl0
,
CAXI4DMAIl0
,
CAXI4DMAl00
,
CAXI4DMAO10
,
CAXI4DMAI10
,
CAXI4DMAl10
,
CAXI4DMAll0
,
CAXI4DMAO00
,
CAXI4DMAI00
,
waitDscrptr
,
waitStrDscrptr
,
CAXI4DMAI1IOI
,
CAXI4DMAlI1l
,
CAXI4DMAOIOOI
,
CAXI4DMAO1IOI
,
CAXI4DMAl0IOI
,
CAXI4DMAI11l
,
CAXI4DMAl11l
,
CAXI4DMAOI
,
CAXI4DMAII
,
CAXI4DMAlI
,
CAXI4DMAOl
,
CAXI4DMAIl
,
CAXI4DMAll
,
CAXI4DMAl0
,
CAXI4DMAO1
,
CAXI4DMAI1
,
CAXI4DMAO0
,
CAXI4DMAI0
,
CAXI4DMAOIlOI
,
CAXI4DMAOOI
,
CAXI4DMAIOI
,
CAXI4DMAIlI
,
CAXI4DMAllI
,
CAXI4DMAO0I
,
CAXI4DMAI0I
,
CAXI4DMAl0I
,
CAXI4DMAO1I
,
CAXI4DMAlOI
,
CAXI4DMAOII
,
CAXI4DMAIII
,
CAXI4DMAlII
,
CAXI4DMAOlI
,
CAXI4DMAI1l1
,
CAXI4DMAl1l1
,
valid
,
CAXI4DMAlIlOI
,
CAXI4DMAOllOI
,
CAXI4DMAIllOI
,
CAXI4DMAlllOI
,
CAXI4DMAO0lOI
,
CAXI4DMAI0lOI
,
CAXI4DMAl0lOI
,
CAXI4DMAO1lOI
,
CAXI4DMAI0IOI
,
CAXI4DMAlll1
,
CAXI4DMAIO01
,
CAXI4DMAII1l
,
CAXI4DMAO1OOI
,
CAXI4DMAOl1l
,
CAXI4DMAIl1l
)
;
parameter
AXI4_STREAM_IF
=
0
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl1OI
=
133
;
parameter
CAXI4DMAl0OI
=
23
;
parameter
NUM_PRI_LVLS
=
1
;
parameter
CAXI4DMAO1OI
=
12
;
parameter
CAXI4DMAI1OI
=
8
;
parameter
PRI_0_NUM_OF_BEATS
=
255
;
parameter
PRI_1_NUM_OF_BEATS
=
127
;
parameter
PRI_2_NUM_OF_BEATS
=
63
;
parameter
PRI_3_NUM_OF_BEATS
=
31
;
parameter
PRI_4_NUM_OF_BEATS
=
15
;
parameter
PRI_5_NUM_OF_BEATS
=
7
;
parameter
PRI_6_NUM_OF_BEATS
=
3
;
parameter
PRI_7_NUM_OF_BEATS
=
0
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAIOlOI
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAlOlOI
;
input
CAXI4DMAI1l
;
input
CAXI4DMAl1l
;
input
CAXI4DMAOO0
;
input
CAXI4DMAIO0
;
input
CAXI4DMAlO0
;
input
CAXI4DMAOI0
;
input
CAXI4DMAII0
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI0
;
input
CAXI4DMAOl0
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIl0
;
input
CAXI4DMAl00
;
input
[
1
:
0
]
CAXI4DMAO10
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAI10
;
input
CAXI4DMAl10
;
input
CAXI4DMAll0
;
input
CAXI4DMAO00
;
input
CAXI4DMAI00
;
input
[
NUM_INT_BDS
-
1
:
0
]
waitDscrptr
;
input
waitStrDscrptr
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAI1IOI
;
input
CAXI4DMAlI1l
;
input
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOIOOI
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
input
CAXI4DMAl0IOI
;
input
CAXI4DMAI11l
;
input
[
31
:
0
]
CAXI4DMAl11l
;
output
CAXI4DMAOI
;
output
CAXI4DMAII
;
output
[
1
:
0
]
CAXI4DMAlI
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOl
;
output
[
31
:
0
]
CAXI4DMAIl
;
output
[
2
:
0
]
CAXI4DMAll
;
output
CAXI4DMAI0
;
output
[
1
:
0
]
CAXI4DMAl0
;
output
[
31
:
0
]
CAXI4DMAO1
;
output
[
2
:
0
]
CAXI4DMAI1
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAO0
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOIlOI
;
output
[
2
:
0
]
CAXI4DMAOOI
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAIOI
;
output
CAXI4DMAIlI
;
output
CAXI4DMAllI
;
output
CAXI4DMAO0I
;
output
[
31
:
0
]
CAXI4DMAI0I
;
output
CAXI4DMAl0I
;
output
[
7
:
0
]
CAXI4DMAO1I
;
output
CAXI4DMAlOI
;
output
[
31
:
0
]
CAXI4DMAOII
;
output
CAXI4DMAIII
;
output
[
31
:
0
]
CAXI4DMAlII
;
output
[
1
:
0
]
CAXI4DMAOlI
;
output
CAXI4DMAI1l1
;
output
CAXI4DMAl1l1
;
output
valid
;
output
CAXI4DMAlIlOI
;
output
CAXI4DMAOllOI
;
output
CAXI4DMAIllOI
;
output
CAXI4DMAlllOI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO0lOI
;
output
CAXI4DMAI0lOI
;
output
[
31
:
0
]
CAXI4DMAl0lOI
;
output
CAXI4DMAO1lOI
;
output
CAXI4DMAI0IOI
;
output
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAlll1
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIO01
;
output
CAXI4DMAII1l
;
output
CAXI4DMAO1OOI
;
output
CAXI4DMAOl1l
;
output
CAXI4DMAIl1l
;
localparam
CAXI4DMAO1llI
=
(
CAXI4DMAl1OI
+
32
+
1
)
;
wire
CAXI4DMAllI0I
;
wire
CAXI4DMAO0I0I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0I0I
;
wire
CAXI4DMAl0IlI
;
wire
CAXI4DMAl0I0I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO1I0I
;
wire
CAXI4DMAI1I0I
;
wire
CAXI4DMAl1I0I
;
wire
CAXI4DMAOOl0I
;
wire
CAXI4DMAIOl0I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlOl0I
;
wire
[
31
:
0
]
CAXI4DMAOIl0I
;
wire
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAIIl0I
;
wire
CAXI4DMAlIl0I
;
wire
CAXI4DMAOll0I
;
wire
CAXI4DMAIll0I
;
wire
CAXI4DMAlll0I
;
wire
CAXI4DMAO0l0I
;
wire
CAXI4DMAI0l0I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl0l0I
;
wire
[
31
:
0
]
CAXI4DMAO1l0I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI1l0I
;
wire
[
31
:
0
]
CAXI4DMAl1l0I
;
wire
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAOO00I
;
wire
CAXI4DMAIO00I
;
wire
CAXI4DMAlO00I
;
wire
CAXI4DMAOI00I
;
wire
CAXI4DMAII00I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlI00I
;
wire
[
31
:
0
]
CAXI4DMAOl00I
;
wire
CAXI4DMAIl00I
;
wire
CAXI4DMAll00I
;
wire
CAXI4DMAO000I
;
wire
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAI000I
;
wire
[
31
:
0
]
CAXI4DMAl000I
;
wire
[
31
:
0
]
CAXI4DMAO100I
;
wire
CAXI4DMAlOllI
;
wire
CAXI4DMAI100I
;
wire
CAXI4DMAlIllI
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOlllI
;
wire
CAXI4DMAIlllI
;
wire
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAl100I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0llI
;
wire
[
CAXI4DMAO1llI
-
1
:
0
]
CAXI4DMAl0llI
;
wire
CAXI4DMAOO10I
;
wire
CAXI4DMAIO10I
;
wire
CAXI4DMAlO10I
;
wire
CAXI4DMAOI10I
;
wire
CAXI4DMAII10I
;
wire
CAXI4DMAlI10I
;
wire
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOl10I
;
wire
[
31
:
0
]
CAXI4DMAIl10I
;
wire
[
7
:
0
]
CAXI4DMAI011
;
wire
CAXI4DMAll10I
;
wire
CAXI4DMAO010I
;
wire
CAXI4DMAI010I
;
wire
CAXI4DMAO0llI
;
wire
CAXI4DMAOIllI
;
wire
CAXI4DMAl010I
;
wire
CAXI4DMAO110I
;
CAXI4DMAI110I
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
)
CAXI4DMAl110I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAlOlOI
(
CAXI4DMAlOlOI
)
,
.CAXI4DMAIOlOI
(
CAXI4DMAIOlOI
)
,
.CAXI4DMAllI0I
(
CAXI4DMAllI0I
)
,
.CAXI4DMAl0IlI
(
CAXI4DMAO0I0I
)
,
.CAXI4DMAI0I0I
(
CAXI4DMAI0I0I
)
)
;
CAXI4DMAOOO1I
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl1OI
(
CAXI4DMAl1OI
)
)
CAXI4DMAIOO1I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAO0I0I
(
CAXI4DMAO0I0I
)
,
.CAXI4DMAlOO1I
(
CAXI4DMAI0I0I
)
,
.CAXI4DMAl0I0I
(
CAXI4DMAl0I0I
)
,
.CAXI4DMAO1I0I
(
CAXI4DMAO1I0I
)
,
.CAXI4DMAI1I0I
(
CAXI4DMAI1I0I
)
,
.CAXI4DMAOIO1I
(
CAXI4DMAlI1l
)
,
.CAXI4DMAIIO1I
(
CAXI4DMAO1IOI
)
,
.CAXI4DMAl0IOI
(
CAXI4DMAl0IOI
)
,
.CAXI4DMAl1I0I
(
CAXI4DMAl1I0I
)
,
.CAXI4DMAOOl0I
(
CAXI4DMAOOl0I
)
,
.CAXI4DMAIOl0I
(
CAXI4DMAIOl0I
)
,
.CAXI4DMAlOl0I
(
CAXI4DMAlOl0I
)
,
.CAXI4DMAOIl0I
(
CAXI4DMAOIl0I
)
,
.CAXI4DMAIIl0I
(
CAXI4DMAIIl0I
)
,
.CAXI4DMAlIl0I
(
CAXI4DMAlIl0I
)
,
.CAXI4DMAllI0I
(
CAXI4DMAllI0I
)
,
.CAXI4DMAOll0I
(
CAXI4DMAOll0I
)
,
.CAXI4DMAIll0I
(
CAXI4DMAIll0I
)
,
.CAXI4DMAI1l0I
(
CAXI4DMAI1l0I
)
,
.CAXI4DMAO010I
(
CAXI4DMAO010I
)
,
.CAXI4DMAI010I
(
CAXI4DMAI010I
)
,
.CAXI4DMAl1l0I
(
CAXI4DMAl1l0I
)
,
.CAXI4DMAl0IlI
(
CAXI4DMAl0IlI
)
,
.CAXI4DMAI1IlI
(
CAXI4DMAlll0I
)
,
.strDscrptr
(
CAXI4DMAO0l0I
)
,
.CAXI4DMAlIO1I
(
CAXI4DMAI0l0I
)
,
.intDscrptrNum
(
CAXI4DMAl0l0I
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAO1l0I
)
,
.CAXI4DMAO1IOI
(
CAXI4DMAOO00I
)
,
.CAXI4DMAOlO1I
(
CAXI4DMAIO00I
)
,
.CAXI4DMAI0IOI
(
CAXI4DMAI0IOI
)
,
.CAXI4DMAIlO1I
(
CAXI4DMAIO01
)
)
;
CAXI4DMAllO1I
#
(
.CAXI4DMAl1OI
(
CAXI4DMAl1OI
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
)
CAXI4DMAO0O1I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAOlO1I
(
CAXI4DMAIO00I
)
,
.CAXI4DMAO1OOI
(
CAXI4DMAI11l
)
,
.CAXI4DMAl11l
(
CAXI4DMAl11l
)
,
.CAXI4DMAI0O1I
(
CAXI4DMAlO00I
)
,
.CAXI4DMAl0O1I
(
CAXI4DMAOI00I
)
,
.CAXI4DMAO1O1I
(
CAXI4DMAII00I
)
,
.CAXI4DMAO1I0I
(
CAXI4DMAlI00I
)
,
.CAXI4DMAI1O1I
(
CAXI4DMAOl00I
)
,
.CAXI4DMAI011
(
CAXI4DMAI011
)
,
.CAXI4DMAI10
(
CAXI4DMAI10
)
,
.CAXI4DMAl10
(
CAXI4DMAl10
)
,
.CAXI4DMAl1O1I
(
CAXI4DMAl00
)
,
.CAXI4DMAO10
(
CAXI4DMAO10
)
,
.CAXI4DMAOOI1I
(
CAXI4DMAII1l
)
,
.CAXI4DMAIOI1I
(
CAXI4DMAO1OOI
)
,
.intDscrptrNum
(
CAXI4DMAlOl0I
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAOIl0I
)
,
.CAXI4DMAO1IOI
(
CAXI4DMAIIl0I
)
,
.CAXI4DMAlI1l
(
CAXI4DMAlIl0I
)
,
.CAXI4DMAI1IlI
(
CAXI4DMAOOl0I
)
,
.CAXI4DMAlOI1I
(
CAXI4DMAIOl0I
)
,
.CAXI4DMAl1I0I
(
CAXI4DMAl1I0I
)
,
.CAXI4DMAl010I
(
CAXI4DMAl010I
)
,
.CAXI4DMAOII1I
(
CAXI4DMAIl00I
)
,
.CAXI4DMAIII1I
(
CAXI4DMAlI10I
)
,
.CAXI4DMAlII1I
(
CAXI4DMAll00I
)
,
.CAXI4DMAOlI1I
(
CAXI4DMAO000I
)
,
.CAXI4DMAIlI
(
CAXI4DMAIlI
)
,
.CAXI4DMAllI
(
CAXI4DMAllI
)
,
.CAXI4DMAO0I
(
CAXI4DMAO0I
)
,
.CAXI4DMAl0I
(
CAXI4DMAl0I
)
,
.CAXI4DMAIlI1I
(
CAXI4DMAI0I
)
,
.CAXI4DMAO1I
(
CAXI4DMAO1I
)
)
;
CAXI4DMAO0IlI
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.NUM_PRI_LVLS
(
NUM_PRI_LVLS
)
,
.CAXI4DMAl1OI
(
CAXI4DMAl1OI
)
,
.CAXI4DMAO1llI
(
CAXI4DMAO1llI
)
,
.AXI4_STREAM_IF
(
AXI4_STREAM_IF
)
)
CAXI4DMAllI1I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAI0IlI
(
CAXI4DMAI1IOI
)
,
.CAXI4DMAOIOOI
(
CAXI4DMAOIOOI
)
,
.CAXI4DMAO1IOI
(
CAXI4DMAOO00I
)
,
.CAXI4DMAl0IlI
(
CAXI4DMAl0IlI
)
,
.CAXI4DMAO1IlI
(
CAXI4DMAO0l0I
)
,
.CAXI4DMAI1IlI
(
CAXI4DMAlll0I
)
,
.CAXI4DMAII0OI
(
CAXI4DMAI0l0I
)
,
.intDscrptrNum
(
CAXI4DMAl0l0I
)
,
.CAXI4DMAl1IlI
(
CAXI4DMAI000I
)
,
.CAXI4DMAOOllI
(
CAXI4DMAl000I
)
,
.CAXI4DMAIOllI
(
CAXI4DMAO100I
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAO1l0I
)
,
.CAXI4DMAlOllI
(
CAXI4DMAlOllI
)
,
.CAXI4DMAOIllI
(
CAXI4DMAOIllI
)
,
.CAXI4DMAIIllI
(
CAXI4DMAI100I
)
,
.CAXI4DMAlIllI
(
CAXI4DMAlIllI
)
,
.CAXI4DMAOlllI
(
CAXI4DMAOlllI
)
,
.waitDscrptr
(
waitDscrptr
)
,
.waitStrDscrptr
(
waitStrDscrptr
)
,
.CAXI4DMAIlllI
(
CAXI4DMAIlllI
)
,
.CAXI4DMAllllI
(
CAXI4DMAl100I
)
,
.CAXI4DMAO0llI
(
CAXI4DMAO0llI
)
,
.CAXI4DMAI0llI
(
CAXI4DMAI0llI
)
,
.CAXI4DMAl0llI
(
CAXI4DMAl0llI
)
,
.CAXI4DMAlll1
(
CAXI4DMAlll1
)
)
;
CAXI4DMAO0I1I
#
(
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
)
CAXI4DMAI0I1I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAIll0I
(
CAXI4DMAIll0I
)
,
.CAXI4DMAl0l0I
(
CAXI4DMAI1l0I
)
,
.CAXI4DMAl0I1I
(
CAXI4DMAO010I
)
,
.CAXI4DMAO0l0I
(
CAXI4DMAI010I
)
,
.CAXI4DMAO1l0I
(
CAXI4DMAl1l0I
)
,
.CAXI4DMAOO10I
(
CAXI4DMAOO10I
)
,
.CAXI4DMAIO10I
(
CAXI4DMAIO10I
)
,
.CAXI4DMAlO10I
(
CAXI4DMAlO10I
)
,
.CAXI4DMAOI10I
(
CAXI4DMAOI10I
)
,
.CAXI4DMAO1I0I
(
CAXI4DMAOl10I
)
,
.CAXI4DMAO1I1I
(
CAXI4DMAll10I
)
,
.CAXI4DMAI1O1I
(
CAXI4DMAIl10I
)
,
.CAXI4DMAOIllI
(
CAXI4DMAO110I
)
,
.valid
(
valid
)
,
.CAXI4DMAlIlOI
(
CAXI4DMAlIlOI
)
,
.CAXI4DMAOllOI
(
CAXI4DMAOllOI
)
,
.CAXI4DMAIllOI
(
CAXI4DMAIllOI
)
,
.CAXI4DMAlllOI
(
CAXI4DMAlllOI
)
,
.intDscrptrNum
(
CAXI4DMAO0lOI
)
,
.CAXI4DMAII0OI
(
CAXI4DMAI0lOI
)
,
.CAXI4DMAlI0OI
(
CAXI4DMAl0lOI
)
,
.strDscrptr
(
CAXI4DMAO1lOI
)
,
.CAXI4DMAI1I1I
(
CAXI4DMAII10I
)
,
.CAXI4DMAI1I0I
(
CAXI4DMAI1I0I
)
)
;
CAXI4DMAl1I1I
#
(
.NUM_INT_BDS
(
NUM_INT_BDS
)
,
.CAXI4DMAOIO1
(
CAXI4DMAOIO1
)
,
.CAXI4DMAl0OI
(
CAXI4DMAl0OI
)
,
.CAXI4DMAO1OI
(
CAXI4DMAO1OI
)
,
.NUM_PRI_LVLS
(
NUM_PRI_LVLS
)
,
.CAXI4DMAI1OI
(
CAXI4DMAI1OI
)
,
.PRI_0_NUM_OF_BEATS
(
PRI_0_NUM_OF_BEATS
)
,
.PRI_1_NUM_OF_BEATS
(
PRI_1_NUM_OF_BEATS
)
,
.PRI_2_NUM_OF_BEATS
(
PRI_2_NUM_OF_BEATS
)
,
.PRI_3_NUM_OF_BEATS
(
PRI_3_NUM_OF_BEATS
)
,
.PRI_4_NUM_OF_BEATS
(
PRI_4_NUM_OF_BEATS
)
,
.PRI_5_NUM_OF_BEATS
(
PRI_5_NUM_OF_BEATS
)
,
.PRI_6_NUM_OF_BEATS
(
PRI_6_NUM_OF_BEATS
)
,
.PRI_7_NUM_OF_BEATS
(
PRI_7_NUM_OF_BEATS
)
,
.AXI4_STREAM_IF
(
AXI4_STREAM_IF
)
)
CAXI4DMAOOl1I
(
.CAXI4DMAI
(
CAXI4DMAI
)
,
.CAXI4DMAl
(
CAXI4DMAl
)
,
.CAXI4DMAIOl1I
(
CAXI4DMAIlllI
)
,
.CAXI4DMAO0llI
(
CAXI4DMAO0llI
)
,
.CAXI4DMAI0llI
(
CAXI4DMAI0llI
)
,
.CAXI4DMAlOl1I
(
CAXI4DMAl0llI
[
165
:
134
]
)
,
.CAXI4DMAOIl1I
(
CAXI4DMAl0llI
[
166
]
)
,
.CAXI4DMAl100I
(
CAXI4DMAl100I
)
,
.CAXI4DMAIIl1I
(
CAXI4DMAl0llI
[
13
]
)
,
.CAXI4DMAlIl1I
(
CAXI4DMAl0llI
[
12
]
)
,
.CAXI4DMAOll1I
(
CAXI4DMAl0llI
[
69
:
38
]
)
,
.CAXI4DMAIll1I
(
CAXI4DMAl0llI
[
1
:
0
]
)
,
.CAXI4DMAlll1I
(
CAXI4DMAl0llI
[
6
:
4
]
)
,
.CAXI4DMAO0l1I
(
CAXI4DMAl0llI
[
37
:
14
]
)
,
.CAXI4DMAI0l1I
(
CAXI4DMAl0llI
[
10
]
)
,
.CAXI4DMAl0l1I
(
CAXI4DMAl0llI
[
11
]
)
,
.CAXI4DMAO1l1I
(
CAXI4DMAl0llI
[
133
:
102
]
)
,
.CAXI4DMAI1l1I
(
CAXI4DMAl0llI
[
101
:
70
]
)
,
.CAXI4DMAl1l1I
(
CAXI4DMAl0llI
[
3
:
2
]
)
,
.CAXI4DMAOO01I
(
CAXI4DMAl0llI
[
9
:
7
]
)
,
.CAXI4DMAII10I
(
CAXI4DMAII10I
)
,
.CAXI4DMAIO01I
(
CAXI4DMAI1l
)
,
.CAXI4DMAlO01I
(
CAXI4DMAl1l
)
,
.CAXI4DMAOI01I
(
CAXI4DMAOO0
)
,
.CAXI4DMAII01I
(
CAXI4DMAIO0
)
,
.CAXI4DMAlO0
(
CAXI4DMAlO0
)
,
.CAXI4DMAOI0
(
CAXI4DMAOI0
)
,
.CAXI4DMAl011
(
CAXI4DMAII0
)
,
.CAXI4DMAO111
(
CAXI4DMAlI0
)
,
.CAXI4DMAOl0
(
CAXI4DMAOl0
)
,
.CAXI4DMAIl0
(
CAXI4DMAIl0
)
,
.CAXI4DMAll0
(
CAXI4DMAll0
)
,
.CAXI4DMAO00
(
CAXI4DMAO00
)
,
.CAXI4DMAI00
(
CAXI4DMAI00
)
,
.CAXI4DMAlI01I
(
CAXI4DMAl010I
)
,
.CAXI4DMAOl01I
(
CAXI4DMAIl00I
)
,
.CAXI4DMAlI10I
(
CAXI4DMAlI10I
)
,
.CAXI4DMAll00I
(
CAXI4DMAll00I
)
,
.CAXI4DMAO000I
(
CAXI4DMAO000I
)
,
.CAXI4DMAIl01I
(
CAXI4DMAOll0I
)
,
.CAXI4DMAlOllI
(
CAXI4DMAlOllI
)
,
.CAXI4DMAOIllI
(
CAXI4DMAOIllI
)
,
.CAXI4DMAIIllI
(
CAXI4DMAI100I
)
,
.CAXI4DMAl1IlI
(
CAXI4DMAI000I
)
,
.CAXI4DMAOOllI
(
CAXI4DMAl000I
)
,
.CAXI4DMAIOllI
(
CAXI4DMAO100I
)
,
.CAXI4DMAIO0lI
(
CAXI4DMAlIllI
)
,
.CAXI4DMAOlllI
(
CAXI4DMAOlllI
)
,
.CAXI4DMAOO10I
(
CAXI4DMAOO10I
)
,
.CAXI4DMAlIlOI
(
CAXI4DMAIO10I
)
,
.CAXI4DMAOllOI
(
CAXI4DMAlO10I
)
,
.CAXI4DMAIllOI
(
CAXI4DMAOI10I
)
,
.CAXI4DMAll01I
(
CAXI4DMAOl10I
)
,
.CAXI4DMAO001I
(
CAXI4DMAll10I
)
,
.CAXI4DMAI001I
(
CAXI4DMAIl10I
)
,
.CAXI4DMAl001I
(
CAXI4DMAO110I
)
,
.CAXI4DMAI1l1
(
CAXI4DMAI1l1
)
,
.CAXI4DMAl1l1
(
CAXI4DMAl1l1
)
,
.CAXI4DMAOI
(
CAXI4DMAOI
)
,
.CAXI4DMAII
(
CAXI4DMAII
)
,
.CAXI4DMAlI
(
CAXI4DMAlI
)
,
.CAXI4DMAOl
(
CAXI4DMAOl
)
,
.CAXI4DMAll
(
CAXI4DMAll
)
,
.CAXI4DMAO101I
(
CAXI4DMAIl
)
,
.CAXI4DMAI0
(
CAXI4DMAI0
)
,
.CAXI4DMAl0
(
CAXI4DMAl0
)
,
.CAXI4DMAI1
(
CAXI4DMAI1
)
,
.CAXI4DMAI101I
(
CAXI4DMAO1
)
,
.CAXI4DMAlOI
(
CAXI4DMAlOI
)
,
.CAXI4DMAOII
(
CAXI4DMAOII
)
,
.CAXI4DMAIII
(
CAXI4DMAIII
)
,
.CAXI4DMAlII
(
CAXI4DMAlII
)
,
.CAXI4DMAOlI
(
CAXI4DMAOlI
)
,
.CAXI4DMAO0
(
CAXI4DMAO0
)
,
.CAXI4DMAOIlOI
(
CAXI4DMAOIlOI
)
,
.CAXI4DMAOOI
(
CAXI4DMAOOI
)
,
.CAXI4DMAIOI
(
CAXI4DMAIOI
)
,
.CAXI4DMAI0O1I
(
CAXI4DMAlO00I
)
,
.CAXI4DMAl0O1I
(
CAXI4DMAOI00I
)
,
.CAXI4DMAO1O1I
(
CAXI4DMAII00I
)
,
.CAXI4DMAlOl0I
(
CAXI4DMAlI00I
)
,
.CAXI4DMAOIl0I
(
CAXI4DMAOl00I
)
,
.CAXI4DMAO1I
(
CAXI4DMAI011
)
,
.CAXI4DMAl0I0I
(
CAXI4DMAl0I0I
)
,
.CAXI4DMAl0l0I
(
CAXI4DMAO1I0I
)
,
.CAXI4DMAOl1l
(
CAXI4DMAOl1l
)
,
.CAXI4DMAIl1l
(
CAXI4DMAIl1l
)
)
;
endmodule
