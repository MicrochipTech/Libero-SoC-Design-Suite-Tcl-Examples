// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAI1lOI
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAll1l
,
CAXI4DMAO01l
,
CAXI4DMAI01l
,
CAXI4DMAl01l
,
CAXI4DMAO11l
,
CAXI4DMAOIO0
,
CAXI4DMAIIO0
,
CAXI4DMAOO0OI
)
;
parameter
CAXI4DMAl110
=
0
;
parameter
CAXI4DMAOOO1
=
0
;
parameter
CAXI4DMAIOO1
=
0
;
parameter
NUM_INT_BDS
=
4
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAll1l
;
input
CAXI4DMAO01l
;
input
[
10
:
0
]
CAXI4DMAI01l
;
input
[
31
:
0
]
CAXI4DMAl01l
;
input
[
3
:
0
]
CAXI4DMAO11l
;
output
[
31
:
0
]
CAXI4DMAOIO0
;
output
CAXI4DMAIIO0
;
output
[
NUM_INT_BDS
-
1
:
0
]
CAXI4DMAOO0OI
;
wire
[
23
:
0
]
CAXI4DMAlIIlI
;
reg
[
31
:
0
]
CAXI4DMAOlIlI
;
localparam
[
10
:
0
]
CAXI4DMAIlIlI
=
11
'h
000
;
localparam
[
10
:
0
]
CAXI4DMAllIlI
=
11
'h
004
;
assign
CAXI4DMAlIIlI
[
7
:
0
]
=
CAXI4DMAIOO1
;
assign
CAXI4DMAlIIlI
[
15
:
8
]
=
CAXI4DMAOOO1
;
assign
CAXI4DMAlIIlI
[
23
:
16
]
=
CAXI4DMAl110
;
assign
CAXI4DMAIIO0
=
1
'b
1
;
assign
CAXI4DMAOIO0
[
31
:
0
]
=
(
CAXI4DMAI01l
==
CAXI4DMAIlIlI
)
?
(
{
{
8
{
1
'b
0
}
}
,
CAXI4DMAlIIlI
[
23
:
0
]
}
)
:
32
'b
0
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOlIlI
<=
32
'b
0
;
end
else
begin
if
(
CAXI4DMAll1l
&
CAXI4DMAO01l
&
(
CAXI4DMAI01l
==
CAXI4DMAllIlI
)
)
begin
if
(
CAXI4DMAO11l
[
0
]
)
begin
CAXI4DMAOlIlI
[
7
:
0
]
<=
CAXI4DMAl01l
[
7
:
0
]
;
end
else
begin
CAXI4DMAOlIlI
[
7
:
0
]
<=
8
'b
0
;
end
if
(
CAXI4DMAO11l
[
1
]
)
begin
CAXI4DMAOlIlI
[
15
:
8
]
<=
CAXI4DMAl01l
[
15
:
8
]
;
end
else
begin
CAXI4DMAOlIlI
[
15
:
8
]
<=
8
'b
0
;
end
if
(
CAXI4DMAO11l
[
2
]
)
begin
CAXI4DMAOlIlI
[
23
:
16
]
<=
CAXI4DMAl01l
[
23
:
16
]
;
end
else
begin
CAXI4DMAOlIlI
[
23
:
16
]
<=
8
'b
0
;
end
if
(
CAXI4DMAO11l
[
3
]
)
begin
CAXI4DMAOlIlI
[
31
:
24
]
<=
CAXI4DMAl01l
[
31
:
24
]
;
end
else
begin
CAXI4DMAOlIlI
[
31
:
24
]
<=
8
'b
0
;
end
end
else
begin
CAXI4DMAOlIlI
<=
32
'b
0
;
end
end
end
assign
CAXI4DMAOO0OI
=
CAXI4DMAOlIlI
;
endmodule
