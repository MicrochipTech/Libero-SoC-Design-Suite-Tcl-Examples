// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAIOIOI
(
CAXI4DMAOIIOI
,
CAXI4DMAIIIOI
,
CAXI4DMAlIIOI
,
CAXI4DMAOlIOI
,
CAXI4DMAIlIOI
,
CAXI4DMAIOI1
,
CAXI4DMAOII1
,
CAXI4DMAlOI1
,
CAXI4DMAlII1
,
CAXI4DMAIII1
,
CAXI4DMAOlI1
,
CAXI4DMAIlI1
,
CAXI4DMAI0OOI
,
CAXI4DMAl0OOI
,
CAXI4DMAll1l
,
CAXI4DMAO01l
,
CAXI4DMAI01l
,
CAXI4DMAl01l
,
CAXI4DMAO11l
,
CAXI4DMAOOIOI
,
CAXI4DMAOIO0
,
CAXI4DMAIIO0
)
;
input
CAXI4DMAOIIOI
;
input
CAXI4DMAIIIOI
;
input
[
10
:
0
]
CAXI4DMAlIIOI
;
input
[
31
:
0
]
CAXI4DMAOlIOI
;
input
[
3
:
0
]
CAXI4DMAIlIOI
;
input
CAXI4DMAIOI1
;
input
[
31
:
0
]
CAXI4DMAOII1
;
input
CAXI4DMAlOI1
;
input
[
31
:
0
]
CAXI4DMAlII1
;
input
CAXI4DMAIII1
;
input
[
31
:
0
]
CAXI4DMAOlI1
;
input
CAXI4DMAIlI1
;
input
[
31
:
0
]
CAXI4DMAI0OOI
;
input
CAXI4DMAl0OOI
;
output
CAXI4DMAll1l
;
output
CAXI4DMAO01l
;
output
[
10
:
0
]
CAXI4DMAI01l
;
output
[
31
:
0
]
CAXI4DMAl01l
;
output
[
3
:
0
]
CAXI4DMAO11l
;
output
CAXI4DMAOOIOI
;
output
[
31
:
0
]
CAXI4DMAOIO0
;
output
CAXI4DMAIIO0
;
assign
CAXI4DMAll1l
=
CAXI4DMAOIIOI
;
assign
CAXI4DMAO01l
=
CAXI4DMAIIIOI
;
assign
CAXI4DMAI01l
=
CAXI4DMAlIIOI
;
assign
CAXI4DMAl01l
=
CAXI4DMAOlIOI
;
assign
CAXI4DMAO11l
=
CAXI4DMAIlIOI
;
assign
CAXI4DMAOIO0
=
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
460
)
?
CAXI4DMAI0OOI
:
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
060
)
?
CAXI4DMAOII1
:
(
CAXI4DMAI01l
[
10
:
0
]
==
11
'h
0
)
?
CAXI4DMAOlI1
:
CAXI4DMAlII1
;
assign
CAXI4DMAIIO0
=
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
460
)
?
CAXI4DMAl0OOI
:
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
060
)
?
CAXI4DMAlOI1
:
(
CAXI4DMAI01l
[
10
:
0
]
==
11
'h
0
)
?
CAXI4DMAIlI1
:
CAXI4DMAIII1
;
assign
CAXI4DMAOOIOI
=
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
460
)
?
1
'b
1
:
(
CAXI4DMAI01l
[
10
:
0
]
>=
11
'h
060
)
?
CAXI4DMAIOI1
:
1
'b
1
;
endmodule
