// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAO
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAOI
,
CAXI4DMAII
,
CAXI4DMAlI
,
CAXI4DMAOl
,
CAXI4DMAIl
,
CAXI4DMAll
,
CAXI4DMAO0
,
CAXI4DMAI0
,
CAXI4DMAl0
,
CAXI4DMAO1
,
CAXI4DMAI1
,
CAXI4DMAl1
,
CAXI4DMAOOI
,
CAXI4DMAIOI
,
CAXI4DMAlOI
,
CAXI4DMAOII
,
CAXI4DMAIII
,
CAXI4DMAlII
,
CAXI4DMAOlI
,
CAXI4DMAIlI
,
CAXI4DMAllI
,
CAXI4DMAO0I
,
CAXI4DMAI0I
,
CAXI4DMAl0I
,
CAXI4DMAO1I
,
CAXI4DMAI1I
,
CAXI4DMAl1I
,
CAXI4DMAOOl
,
CAXI4DMAIOl
,
CAXI4DMAlOl
,
CAXI4DMAOIl
,
CAXI4DMAIIl
,
CAXI4DMAlIl
,
CAXI4DMAOll
,
CAXI4DMAIll
,
CAXI4DMAlll
,
CAXI4DMAO0l
,
CAXI4DMAI0l
,
CAXI4DMAl0l
,
CAXI4DMAO1l
,
CAXI4DMAI1l
,
CAXI4DMAl1l
,
CAXI4DMAOO0
,
CAXI4DMAIO0
,
CAXI4DMAlO0
,
CAXI4DMAOI0
,
CAXI4DMAII0
,
CAXI4DMAlI0
,
CAXI4DMAOl0
,
CAXI4DMAIl0
,
CAXI4DMAll0
,
CAXI4DMAO00
,
CAXI4DMAI00
,
CAXI4DMAl00
,
CAXI4DMAO10
,
CAXI4DMAI10
,
CAXI4DMAl10
,
CAXI4DMAOO1
,
CAXI4DMAIO1
,
CAXI4DMAlO1
,
CAXI4DMAOI1
,
CAXI4DMAII1
,
CAXI4DMAlI1
,
CAXI4DMAOl1
,
CAXI4DMAIl1
,
CAXI4DMAll1
,
CAXI4DMAO01
,
CAXI4DMAI01
,
CAXI4DMAl01
,
CAXI4DMAO11
,
CAXI4DMAI11
,
CAXI4DMAl11
,
CAXI4DMAOOOI
,
CAXI4DMAIOOI
,
CAXI4DMAlOOI
,
CAXI4DMAOIOI
,
CAXI4DMAIIOI
,
CAXI4DMAlIOI
,
CAXI4DMAOlOI
,
CAXI4DMAIlOI
,
CAXI4DMAllOI
,
CAXI4DMAO0OI
,
CAXI4DMAI0OI
)
;
parameter
AXI4_STREAM_IF
=
0
;
parameter
AXI_DMA_DWIDTH
=
0
;
parameter
CAXI4DMAl0OI
=
23
;
parameter
CAXI4DMAO1OI
=
12
;
parameter
CAXI4DMAI1OI
=
8
;
parameter
CAXI4DMAl1OI
=
160
;
parameter
CAXI4DMAOOII
=
256
;
parameter
ID_WIDTH
=
1
;
function
integer
CAXI4DMAIOII
;
input
integer
CAXI4DMAlOII
;
integer
CAXI4DMAOIII
,
CAXI4DMAIIII
,
CAXI4DMAlIII
;
begin
CAXI4DMAIIII
=
1
;
CAXI4DMAlIII
=
0
;
CAXI4DMAOIII
=
CAXI4DMAlOII
+
1
;
while
(
CAXI4DMAIIII
<
CAXI4DMAOIII
)
begin
CAXI4DMAIIII
=
CAXI4DMAIIII
*
2
;
CAXI4DMAlIII
=
CAXI4DMAlIII
+
1
;
end
CAXI4DMAIOII
=
CAXI4DMAlIII
;
end
endfunction
localparam
CAXI4DMAOlII
=
CAXI4DMAIOII
(
AXI_DMA_DWIDTH
/
8
)
;
localparam
CAXI4DMAIlII
=
CAXI4DMAIOII
(
(
AXI_DMA_DWIDTH
/
8
)
-
1
)
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAOI
;
input
CAXI4DMAII
;
input
[
1
:
0
]
CAXI4DMAlI
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOl
;
input
[
31
:
0
]
CAXI4DMAIl
;
input
[
2
:
0
]
CAXI4DMAll
;
input
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAO0
;
input
CAXI4DMAI0
;
input
[
1
:
0
]
CAXI4DMAl0
;
input
[
31
:
0
]
CAXI4DMAO1
;
input
[
2
:
0
]
CAXI4DMAI1
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl1
;
input
[
2
:
0
]
CAXI4DMAOOI
;
input
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAIOI
;
input
CAXI4DMAlOI
;
input
[
31
:
0
]
CAXI4DMAOII
;
input
CAXI4DMAIII
;
input
[
31
:
0
]
CAXI4DMAlII
;
input
[
1
:
0
]
CAXI4DMAOlI
;
input
CAXI4DMAIlI
;
input
CAXI4DMAllI
;
input
CAXI4DMAO0I
;
input
[
31
:
0
]
CAXI4DMAI0I
;
input
CAXI4DMAl0I
;
input
[
7
:
0
]
CAXI4DMAO1I
;
input
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAI1I
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAl1I
;
input
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAOOl
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIOl
;
input
[
1
:
0
]
CAXI4DMAlOl
;
input
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAOIl
;
input
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAIIl
;
input
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAlIl
;
input
CAXI4DMAOll
;
input
CAXI4DMAIll
;
input
CAXI4DMAlll
;
input
CAXI4DMAO0l
;
input
CAXI4DMAI0l
;
input
[
1
:
0
]
CAXI4DMAl0l
;
input
CAXI4DMAO1l
;
output
CAXI4DMAI1l
;
output
CAXI4DMAl1l
;
output
CAXI4DMAOO0
;
output
CAXI4DMAIO0
;
output
CAXI4DMAlO0
;
output
CAXI4DMAOI0
;
output
CAXI4DMAII0
;
output
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI0
;
output
CAXI4DMAOl0
;
output
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIl0
;
output
reg
CAXI4DMAll0
;
output
reg
CAXI4DMAO00
;
output
reg
CAXI4DMAI00
;
output
reg
CAXI4DMAl00
;
output
reg
[
1
:
0
]
CAXI4DMAO10
;
output
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAI10
;
output
reg
CAXI4DMAl10
;
output
CAXI4DMAOO1
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAIO1
;
output
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAlO1
;
output
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAOI1
;
output
reg
CAXI4DMAII1
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAlI1
;
output
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAOl1
;
output
reg
CAXI4DMAIl1
;
output
CAXI4DMAll1
;
output
CAXI4DMAO01
;
output
CAXI4DMAI01
;
output
CAXI4DMAl01
;
output
CAXI4DMAO11
;
output
CAXI4DMAI11
;
output
[
31
:
0
]
CAXI4DMAl11
;
output
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAOOOI
;
output
[
7
:
0
]
CAXI4DMAIOOI
;
output
[
2
:
0
]
CAXI4DMAlOOI
;
output
[
1
:
0
]
CAXI4DMAOIOI
;
output
[
(
AXI_DMA_DWIDTH
/
8
)
-
1
:
0
]
CAXI4DMAIIOI
;
output
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAlIOI
;
output
[
31
:
0
]
CAXI4DMAOlOI
;
output
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAIlOI
;
output
[
7
:
0
]
CAXI4DMAllOI
;
output
[
2
:
0
]
CAXI4DMAO0OI
;
output
[
1
:
0
]
CAXI4DMAI0OI
;
reg
[
12
:
0
]
CAXI4DMAllII
;
reg
[
12
:
0
]
CAXI4DMAO0II
;
reg
[
12
:
0
]
CAXI4DMAI0II
;
reg
[
12
:
0
]
CAXI4DMAl0II
;
wire
[
7
:
0
]
CAXI4DMAO1II
;
reg
CAXI4DMAI1II
;
reg
CAXI4DMAl1II
;
reg
[
31
:
0
]
CAXI4DMAOOlI
;
reg
[
31
:
0
]
CAXI4DMAIOlI
;
reg
[
2
:
0
]
CAXI4DMAlOlI
;
reg
[
2
:
0
]
CAXI4DMAOIlI
;
reg
[
1
:
0
]
CAXI4DMAIIlI
;
reg
[
1
:
0
]
CAXI4DMAlIlI
;
reg
[
7
:
0
]
CAXI4DMAOllI
;
reg
[
7
:
0
]
CAXI4DMAIllI
;
reg
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAlllI
;
reg
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAO0lI
;
reg
CAXI4DMAI0lI
;
reg
CAXI4DMAl0lI
;
reg
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAO1lI
;
reg
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAI1lI
;
reg
CAXI4DMAl1lI
;
reg
CAXI4DMAOO0I
;
reg
[
(
AXI_DMA_DWIDTH
/
8
)
-
1
:
0
]
CAXI4DMAIO0I
;
reg
[
(
AXI_DMA_DWIDTH
/
8
)
-
1
:
0
]
CAXI4DMAlO0I
;
reg
CAXI4DMAOI0I
;
reg
CAXI4DMAII0I
;
reg
CAXI4DMAlO0
;
reg
CAXI4DMAOI0
;
reg
CAXI4DMAI1l
;
reg
CAXI4DMAOO0
;
reg
[
7
:
0
]
CAXI4DMAlI0I
;
reg
[
7
:
0
]
CAXI4DMAOl0I
;
reg
[
8
:
0
]
CAXI4DMAIl0I
;
reg
[
8
:
0
]
CAXI4DMAll0I
;
reg
[
7
:
0
]
CAXI4DMAO00I
;
reg
[
7
:
0
]
CAXI4DMAI00I
;
reg
CAXI4DMAl00I
;
reg
CAXI4DMAO10I
;
reg
[
31
:
0
]
CAXI4DMAI10I
;
reg
[
31
:
0
]
CAXI4DMAl10I
;
reg
[
2
:
0
]
CAXI4DMAOO1I
;
reg
[
2
:
0
]
CAXI4DMAIO1I
;
reg
[
1
:
0
]
CAXI4DMAlO1I
;
reg
[
1
:
0
]
CAXI4DMAOI1I
;
reg
[
7
:
0
]
CAXI4DMAII1I
;
reg
[
7
:
0
]
CAXI4DMAlI1I
;
reg
CAXI4DMAOl1I
;
reg
CAXI4DMAIl1I
;
reg
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI0
;
reg
CAXI4DMAII0
;
reg
[
7
:
0
]
CAXI4DMAll1I
;
reg
[
7
:
0
]
CAXI4DMAO01I
;
reg
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAI01I
;
reg
[
ID_WIDTH
-
1
:
0
]
CAXI4DMAl01I
;
reg
CAXI4DMAl1l
;
reg
CAXI4DMAIO0
;
reg
[
7
:
0
]
CAXI4DMAO11I
;
reg
[
7
:
0
]
CAXI4DMAI11I
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAl11I
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOOOl
;
reg
[
31
:
0
]
CAXI4DMAIOOl
;
reg
[
31
:
0
]
CAXI4DMAlOOl
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOIOl
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIIOl
;
reg
[
1
:
0
]
CAXI4DMAlIOl
;
reg
[
1
:
0
]
CAXI4DMAOlOl
;
reg
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIlOl
;
reg
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAllOl
;
reg
CAXI4DMAO0Ol
;
reg
CAXI4DMAI0Ol
;
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAl0Ol
;
reg
CAXI4DMAO1Ol
;
reg
[
1
:
0
]
CAXI4DMAI1Ol
;
reg
CAXI4DMAl1Ol
;
reg
CAXI4DMAOOIl
;
reg
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAIOIl
;
reg
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAlOIl
;
reg
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAOIIl
;
reg
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAIIIl
;
reg
CAXI4DMAlIIl
;
reg
CAXI4DMAOlIl
;
reg
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAIlIl
;
reg
[
CAXI4DMAOlII
-
1
:
0
]
CAXI4DMAllIl
;
reg
[
1
:
0
]
CAXI4DMAO0Il
;
reg
[
1
:
0
]
CAXI4DMAI0Il
;
reg
CAXI4DMAl0Il
;
reg
CAXI4DMAO1Il
;
reg
[
AXI_DMA_DWIDTH
-
1
:
0
]
CAXI4DMAI1Il
;
reg
CAXI4DMAl1Il
;
reg
CAXI4DMAOOll
;
reg
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAIOll
;
reg
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlOll
;
reg
CAXI4DMAOIll
;
reg
CAXI4DMAIIll
;
localparam
[
12
:
0
]
CAXI4DMAlIll
=
13
'b
0000000000001
;
localparam
[
12
:
0
]
CAXI4DMAOlll
=
13
'b
0000000000010
;
localparam
[
12
:
0
]
CAXI4DMAIlll
=
13
'b
0000000000100
;
localparam
[
12
:
0
]
CAXI4DMAllll
=
13
'b
0000000001000
;
localparam
[
12
:
0
]
CAXI4DMAO0ll
=
13
'b
0000000010000
;
localparam
[
12
:
0
]
CAXI4DMAI0ll
=
13
'b
0000000100000
;
localparam
[
12
:
0
]
CAXI4DMAl0ll
=
13
'b
0000001000000
;
localparam
[
12
:
0
]
CAXI4DMAO1ll
=
13
'b
0000010000000
;
localparam
[
12
:
0
]
CAXI4DMAI1ll
=
13
'b
0000100000000
;
localparam
[
12
:
0
]
CAXI4DMAl1ll
=
13
'b
0001000000000
;
localparam
[
12
:
0
]
CAXI4DMAOO0l
=
13
'b
0010000000000
;
localparam
[
12
:
0
]
CAXI4DMAIO0l
=
13
'b
0100000000000
;
localparam
[
12
:
0
]
CAXI4DMAlO0l
=
13
'b
1000000000000
;
localparam
[
12
:
0
]
CAXI4DMAOI0l
=
13
'b
0000000000001
;
localparam
[
12
:
0
]
CAXI4DMAII0l
=
13
'b
0000000000010
;
localparam
[
12
:
0
]
CAXI4DMAlI0l
=
13
'b
0000000000100
;
localparam
[
12
:
0
]
CAXI4DMAOl0l
=
13
'b
0000000001000
;
localparam
[
12
:
0
]
CAXI4DMAIl0l
=
13
'b
0000000010000
;
localparam
[
12
:
0
]
CAXI4DMAll0l
=
13
'b
0000000100000
;
localparam
[
12
:
0
]
CAXI4DMAO00l
=
13
'b
0000001000000
;
localparam
[
12
:
0
]
CAXI4DMAI00l
=
13
'b
0000010000000
;
localparam
[
12
:
0
]
CAXI4DMAl00l
=
13
'b
0000100000000
;
localparam
[
12
:
0
]
CAXI4DMAO10l
=
13
'b
0001000000000
;
localparam
[
12
:
0
]
CAXI4DMAI10l
=
13
'b
0010000000000
;
localparam
[
12
:
0
]
CAXI4DMAl10l
=
13
'b
0100000000000
;
localparam
[
12
:
0
]
CAXI4DMAOO1l
=
13
'b
1000000000000
;
generate
if
(
AXI_DMA_DWIDTH
==
32
)
begin
assign
CAXI4DMAO1II
=
(
(
CAXI4DMAOIOl
[
1
:
0
]
)
==
1
)
?
4
'b
0001
:
(
(
CAXI4DMAOIOl
[
1
:
0
]
)
==
2
)
?
4
'b
0011
:
(
(
CAXI4DMAOIOl
[
1
:
0
]
)
==
3
)
?
4
'b
0111
:
4
'b
1111
;
end
else
if
(
AXI_DMA_DWIDTH
==
64
)
begin
assign
CAXI4DMAO1II
=
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
1
)
?
8
'b
0000_0001
:
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
2
)
?
8
'b
0000_0011
:
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
3
)
?
8
'b
0000_0111
:
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
4
)
?
8
'b
0000_1111
:
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
5
)
?
8
'b
0001_1111
:
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
6
)
?
8
'b
0011_1111
:
(
(
CAXI4DMAOIOl
[
2
:
0
]
)
==
7
)
?
8
'b
0111_1111
:
8
'b
1111_1111
;
end
else
if
(
AXI_DMA_DWIDTH
==
128
)
begin
assign
CAXI4DMAO1II
=
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
1
)
?
16
'b
0000_0000_0000_0001
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
2
)
?
16
'b
0000_0000_0000_0011
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
3
)
?
16
'b
0000_0000_0000_0111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
4
)
?
16
'b
0000_0000_0000_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
5
)
?
16
'b
0000_0000_0001_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
6
)
?
16
'b
0000_0000_0011_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
7
)
?
16
'b
0000_0000_0111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
8
)
?
16
'b
0000_0000_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
9
)
?
16
'b
0000_0001_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
10
)
?
16
'b
0000_0011_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
11
)
?
16
'b
0000_0111_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
12
)
?
16
'b
0000_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
13
)
?
16
'b
0001_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
14
)
?
16
'b
0011_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
3
:
0
]
)
==
15
)
?
16
'b
0111_1111_1111_1111
:
16
'b
1111_1111_1111_1111
;
end
else
if
(
AXI_DMA_DWIDTH
==
256
)
begin
assign
CAXI4DMAO1II
=
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
1
)
?
32
'b
0000_0000_0000_0000_0000_0000_0000_0001
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
2
)
?
32
'b
0000_0000_0000_0000_0000_0000_0000_0011
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
3
)
?
32
'b
0000_0000_0000_0000_0000_0000_0000_0111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
4
)
?
32
'b
0000_0000_0000_0000_0000_0000_0000_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
5
)
?
32
'b
0000_0000_0000_0000_0000_0000_0001_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
6
)
?
32
'b
0000_0000_0000_0000_0000_0000_0011_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
7
)
?
32
'b
0000_0000_0000_0000_0000_0000_0111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
8
)
?
32
'b
0000_0000_0000_0000_0000_0000_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
9
)
?
32
'b
0000_0000_0000_0000_0000_0001_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
10
)
?
32
'b
0000_0000_0000_0000_0000_0011_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
11
)
?
32
'b
0000_0000_0000_0000_0000_0111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
12
)
?
32
'b
0000_0000_0000_0000_0000_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
13
)
?
32
'b
0000_0000_0000_0000_0001_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
14
)
?
32
'b
0000_0000_0000_0000_0011_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
15
)
?
32
'b
0000_0000_0000_0000_0111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
16
)
?
32
'b
0000_0000_0000_0000_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
17
)
?
32
'b
0000_0000_0000_0001_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
18
)
?
32
'b
0000_0000_0000_0011_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
19
)
?
32
'b
0000_0000_0000_0111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
20
)
?
32
'b
0000_0000_0000_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
21
)
?
32
'b
0000_0000_0001_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
22
)
?
32
'b
0000_0000_0011_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
23
)
?
32
'b
0000_0000_0111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
24
)
?
32
'b
0000_0000_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
25
)
?
32
'b
0000_0001_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
26
)
?
32
'b
0000_0011_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
27
)
?
32
'b
0000_0111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
28
)
?
32
'b
0000_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
29
)
?
32
'b
0001_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
30
)
?
32
'b
0011_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
4
:
0
]
)
==
31
)
?
32
'b
0111_1111_1111_1111_1111_1111_1111_1111
:
32
'b
1111_1111_1111_1111_1111_1111_1111_1111
;
end
else
if
(
AXI_DMA_DWIDTH
==
512
)
begin
assign
CAXI4DMAO1II
=
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
1
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
2
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
3
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
4
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
5
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
6
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
7
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
8
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
9
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
10
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
11
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
12
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
13
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
14
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
15
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
16
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
17
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
18
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
19
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
20
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
21
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
22
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
23
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
24
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
25
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
26
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
27
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
28
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
29
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
30
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
31
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
32
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
33
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
34
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
35
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
36
)
?
64
'b
0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
37
)
?
64
'b
0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
38
)
?
64
'b
0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
39
)
?
64
'b
0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
40
)
?
64
'b
0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
41
)
?
64
'b
0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
42
)
?
64
'b
0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
43
)
?
64
'b
0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
44
)
?
64
'b
0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
45
)
?
64
'b
0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
46
)
?
64
'b
0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
47
)
?
64
'b
0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
48
)
?
64
'b
0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
49
)
?
64
'b
0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
50
)
?
64
'b
0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
51
)
?
64
'b
0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
52
)
?
64
'b
0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
53
)
?
64
'b
0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
54
)
?
64
'b
0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
55
)
?
64
'b
0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
56
)
?
64
'b
0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
57
)
?
64
'b
0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
58
)
?
64
'b
0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
59
)
?
64
'b
0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
60
)
?
64
'b
0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
61
)
?
64
'b
0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
62
)
?
64
'b
0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
(
(
CAXI4DMAOIOl
[
5
:
0
]
)
==
63
)
?
64
'b
0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
:
64
'b
1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111
;
end
endgenerate
always
@
(
*
)
begin
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAl0Il
==
1
'b
1
)
)
begin
CAXI4DMAI1Il
=
CAXI4DMAOOl
;
CAXI4DMAIl1
=
CAXI4DMAlIIl
;
CAXI4DMAII1
=
1
'b
0
;
end
else
begin
CAXI4DMAI1Il
=
CAXI4DMAI1I
;
CAXI4DMAII1
=
CAXI4DMAlIIl
;
CAXI4DMAIl1
=
1
'b
0
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI0II
<=
CAXI4DMAOI0l
;
end
else
begin
CAXI4DMAI0II
<=
CAXI4DMAl0II
;
end
end
always
@
(
*
)
begin
CAXI4DMAl1II
=
1
'b
0
;
CAXI4DMAIOlI
=
CAXI4DMAOOlI
;
CAXI4DMAO0lI
=
{
ID_WIDTH
{
1
'b
0
}
}
;
CAXI4DMAIllI
=
CAXI4DMAOllI
;
CAXI4DMAOIlI
=
CAXI4DMAlOlI
;
CAXI4DMAlIlI
=
CAXI4DMAIIlI
;
CAXI4DMAl0lI
=
1
'b
0
;
CAXI4DMAlO0I
=
CAXI4DMAIO0I
;
CAXI4DMAI1lI
=
CAXI4DMAO1lI
;
CAXI4DMAOO0I
=
CAXI4DMAl1lI
;
CAXI4DMAII0I
=
1
'b
0
;
CAXI4DMAOlIl
=
1
'b
0
;
CAXI4DMAI00I
=
CAXI4DMAO00I
;
CAXI4DMAllIl
=
{
CAXI4DMAOlII
{
1
'b
0
}
}
;
CAXI4DMAll0I
=
CAXI4DMAIl0I
;
CAXI4DMAlO0
=
1
'b
0
;
CAXI4DMAI1l
=
1
'b
0
;
CAXI4DMAOI0
=
1
'b
0
;
CAXI4DMAOO0
=
1
'b
0
;
CAXI4DMAOl0I
=
CAXI4DMAlI0I
;
CAXI4DMAlOOl
=
CAXI4DMAIOOl
;
CAXI4DMAIIOl
=
CAXI4DMAOIOl
;
CAXI4DMAOlOl
=
CAXI4DMAlIOl
;
CAXI4DMAllOl
=
CAXI4DMAIlOl
;
CAXI4DMAO0Ol
=
1
'b
0
;
CAXI4DMAO1Il
=
CAXI4DMAl0Il
;
CAXI4DMAOOll
=
1
'b
0
;
CAXI4DMAlOll
=
CAXI4DMAIOll
;
CAXI4DMAI00
=
1
'b
0
;
case
(
CAXI4DMAI0II
)
CAXI4DMAOI0l
:
begin
if
(
CAXI4DMAOI
)
begin
CAXI4DMAO1Il
=
CAXI4DMAI0
;
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAI0
==
1
'b
1
)
)
begin
CAXI4DMAIIOl
=
CAXI4DMAl1
;
CAXI4DMAlOOl
=
CAXI4DMAO1
;
if
(
CAXI4DMAl0
==
2
'b
10
)
begin
CAXI4DMAOlOl
=
2
'b
00
;
end
else
begin
CAXI4DMAOlOl
=
2
'b
01
;
end
if
(
(
CAXI4DMAl1
>=
(
1
+
(
CAXI4DMAIOI
<<
CAXI4DMAIlII
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
(
1
+
CAXI4DMAIOI
)
<<
CAXI4DMAIlII
)
)
)
begin
CAXI4DMAOl0I
=
CAXI4DMAIOI
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
127
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
128
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
127
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
63
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
64
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
63
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
31
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
32
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
31
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
15
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
16
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
15
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
7
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
8
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
7
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
3
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
4
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
3
;
end
else
begin
CAXI4DMAOl0I
=
8
'd
0
;
end
CAXI4DMAOOll
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAOO1l
;
end
else
begin
CAXI4DMAIIOl
=
CAXI4DMAl1
;
CAXI4DMAlOOl
=
CAXI4DMAO1
;
if
(
CAXI4DMAl1I
>=
CAXI4DMAl1
)
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAIOlI
=
CAXI4DMAO1
;
CAXI4DMAOIlI
=
CAXI4DMAIlII
;
if
(
CAXI4DMAl0
==
2
'b
10
)
begin
CAXI4DMAlIlI
=
2
'b
00
;
end
else
begin
CAXI4DMAlIlI
=
2
'b
01
;
end
if
(
(
CAXI4DMAl1
>=
(
1
+
(
CAXI4DMAIOI
<<
CAXI4DMAIlII
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
(
1
+
CAXI4DMAIOI
)
<<
CAXI4DMAIlII
)
)
)
begin
CAXI4DMAIllI
=
CAXI4DMAIOI
;
CAXI4DMAOl0I
=
CAXI4DMAIOI
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
127
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
128
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAIllI
=
8
'd
127
;
CAXI4DMAOl0I
=
8
'd
127
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
63
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
64
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAIllI
=
8
'd
63
;
CAXI4DMAOl0I
=
8
'd
63
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
31
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
32
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAIllI
=
8
'd
31
;
CAXI4DMAOl0I
=
8
'd
31
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
15
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
16
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAIllI
=
8
'd
15
;
CAXI4DMAOl0I
=
8
'd
15
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
7
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
8
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAIllI
=
8
'd
7
;
CAXI4DMAOl0I
=
8
'd
7
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
3
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
4
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAIllI
=
8
'd
3
;
CAXI4DMAOl0I
=
8
'd
3
;
end
else
begin
CAXI4DMAIllI
=
8
'd
0
;
CAXI4DMAOl0I
=
8
'd
0
;
end
CAXI4DMAl0II
=
CAXI4DMAII0l
;
end
else
begin
if
(
CAXI4DMAl0
==
2
'b
10
)
begin
CAXI4DMAOlOl
=
2
'b
00
;
end
else
begin
CAXI4DMAOlOl
=
2
'b
01
;
end
if
(
(
CAXI4DMAl1
>=
(
1
+
(
CAXI4DMAIOI
<<
CAXI4DMAIlII
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
(
1
+
CAXI4DMAIOI
)
<<
CAXI4DMAIlII
)
)
)
begin
CAXI4DMAOl0I
=
CAXI4DMAIOI
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
127
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
128
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
127
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
63
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
64
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
63
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
31
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
32
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
31
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
15
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
16
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
15
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
7
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
8
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
7
;
end
else
if
(
(
CAXI4DMAl1
>=
(
1
+
(
3
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAO1
[
11
:
0
]
<=
13
'd
4096
-
(
4
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
3
;
end
else
begin
CAXI4DMAOl0I
=
8
'd
0
;
end
CAXI4DMAl0II
=
CAXI4DMAlI0l
;
end
end
end
else
if
(
CAXI4DMAl0I
)
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAIOlI
=
CAXI4DMAI0I
;
CAXI4DMAOIlI
=
CAXI4DMAIlII
;
CAXI4DMAlIlI
=
2
'b
01
;
CAXI4DMAIllI
=
8
'd
0
;
CAXI4DMAl0II
=
CAXI4DMAO00l
;
end
else
if
(
CAXI4DMAIII
)
begin
CAXI4DMAIOlI
=
CAXI4DMAlII
;
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAOIlI
=
CAXI4DMAIlII
;
CAXI4DMAlIlI
=
2
'b
01
;
CAXI4DMAIllI
=
8
'd
0
;
CAXI4DMAO1Il
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAO00l
;
end
else
begin
CAXI4DMAl0II
=
CAXI4DMAOI0l
;
end
end
CAXI4DMAlI0l
:
begin
if
(
CAXI4DMAl1I
>=
CAXI4DMAOIOl
)
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAIOlI
=
CAXI4DMAIOOl
;
CAXI4DMAOIlI
=
CAXI4DMAIlII
;
CAXI4DMAIllI
=
CAXI4DMAlI0I
;
CAXI4DMAlIlI
=
CAXI4DMAlIOl
;
CAXI4DMAl0II
=
CAXI4DMAII0l
;
end
else
begin
CAXI4DMAl0II
=
CAXI4DMAlI0l
;
end
end
CAXI4DMAII0l
:
begin
if
(
CAXI4DMAll1
&
CAXI4DMAOll
)
begin
CAXI4DMAIOlI
=
32
'b
0
;
CAXI4DMAIllI
=
8
'b
0
;
CAXI4DMAOIlI
=
3
'b
0
;
CAXI4DMAlIlI
=
2
'b
0
;
CAXI4DMAI1lI
=
CAXI4DMAI1Il
;
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAOlIl
=
1
'b
1
;
if
(
CAXI4DMAIl0I
==
CAXI4DMAlI0I
)
begin
CAXI4DMAOO0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAI10l
;
if
(
(
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
!=
{
CAXI4DMAIlII
{
1
'b
0
}
}
)
&&
(
CAXI4DMAOIOl
<=
(
AXI_DMA_DWIDTH
/
8
)
)
)
begin
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
;
CAXI4DMAllIl
=
{
1
'b
0
,
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
}
;
CAXI4DMAlO0I
=
CAXI4DMAO1II
;
end
else
begin
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAllIl
=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
1
}
}
;
end
end
else
begin
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAI00I
=
CAXI4DMAO00I
+
1
'b
1
;
CAXI4DMAllIl
=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
1
}
}
;
if
(
CAXI4DMAIl0I
==
CAXI4DMAlI0I
-
1
)
begin
CAXI4DMAl0II
=
CAXI4DMAO10l
;
end
else
begin
CAXI4DMAl0II
=
CAXI4DMAOl0l
;
end
end
end
else
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAII0l
;
end
end
CAXI4DMAOl0l
:
begin
if
(
CAXI4DMAO01
&
CAXI4DMAIll
)
begin
CAXI4DMAll0I
=
CAXI4DMAIl0I
+
1
'b
1
;
CAXI4DMAI1lI
=
CAXI4DMAI1Il
;
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAOlIl
=
1
'b
1
;
CAXI4DMAI00I
=
CAXI4DMAO00I
+
1
'b
1
;
CAXI4DMAllIl
=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
1
}
}
;
if
(
CAXI4DMAIl0I
==
CAXI4DMAlI0I
-
2
'd
2
)
begin
CAXI4DMAl0II
=
CAXI4DMAO10l
;
end
else
begin
CAXI4DMAl0II
=
CAXI4DMAOl0l
;
end
end
else
begin
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAOl0l
;
end
end
CAXI4DMAO10l
:
begin
if
(
CAXI4DMAO01
&
CAXI4DMAIll
)
begin
CAXI4DMAll0I
=
CAXI4DMAIl0I
+
1
'b
1
;
CAXI4DMAI1lI
=
CAXI4DMAI1Il
;
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAOlIl
=
1
'b
1
;
CAXI4DMAOO0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAI10l
;
if
(
CAXI4DMAOIOl
<=
(
CAXI4DMAIlOl
+
(
AXI_DMA_DWIDTH
/
8
)
)
)
begin
if
(
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
==
{
CAXI4DMAIlII
{
1
'b
0
}
}
)
begin
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAllIl
=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
1
}
}
;
end
else
begin
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
;
CAXI4DMAllIl
=
{
1
'b
0
,
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
}
;
CAXI4DMAlO0I
=
CAXI4DMAO1II
;
end
end
else
begin
CAXI4DMAllOl
=
CAXI4DMAIlOl
+
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAllIl
=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
1
}
}
;
end
end
else
begin
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAO10l
;
end
end
CAXI4DMAI10l
:
begin
if
(
CAXI4DMAO01
&
CAXI4DMAIll
)
begin
CAXI4DMAll0I
=
9
'b
0
;
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
0
}
}
;
CAXI4DMAI1lI
=
{
AXI_DMA_DWIDTH
{
1
'b
0
}
}
;
CAXI4DMAOO0I
=
1
'b
0
;
CAXI4DMAII0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAIl0l
;
end
else
begin
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAI10l
;
end
end
CAXI4DMAIl0l
:
begin
if
(
CAXI4DMAlll
&
CAXI4DMAl01
)
begin
if
(
CAXI4DMAlOl
==
2
'b
00
)
begin
if
(
CAXI4DMAOIOl
==
CAXI4DMAIlOl
)
begin
CAXI4DMAI00I
=
8
'b
0
;
CAXI4DMAllOl
=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
CAXI4DMAl0II
=
CAXI4DMAOI0l
;
if
(
(
CAXI4DMAl0Il
==
1
'b
1
)
&&
(
AXI4_STREAM_IF
==
1
)
)
begin
CAXI4DMAlO0
=
1
'b
1
;
CAXI4DMAO1Il
=
1
'b
0
;
end
else
begin
CAXI4DMAI1l
=
1
'b
1
;
end
end
else
begin
CAXI4DMAI00I
=
CAXI4DMAO00I
+
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAll0l
;
end
end
else
begin
CAXI4DMAI00I
=
8
'b
0
;
CAXI4DMAllOl
=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
CAXI4DMAl0II
=
CAXI4DMAOI0l
;
if
(
(
CAXI4DMAl0Il
==
1
'b
1
)
&&
(
AXI4_STREAM_IF
==
1
)
)
begin
CAXI4DMAOI0
=
1
'b
1
;
CAXI4DMAO1Il
=
1
'b
0
;
end
else
begin
CAXI4DMAOO0
=
1
'b
1
;
end
end
end
else
begin
CAXI4DMAII0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAIl0l
;
end
end
CAXI4DMAll0l
:
begin
CAXI4DMAllOl
=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
CAXI4DMAIIOl
=
CAXI4DMAOIOl
-
CAXI4DMAIlOl
;
if
(
CAXI4DMAl0
==
2
'b
10
)
begin
end
else
begin
CAXI4DMAIOlI
=
CAXI4DMAIOOl
+
CAXI4DMAIlOl
;
CAXI4DMAlOOl
=
CAXI4DMAIOOl
+
CAXI4DMAIlOl
;
end
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
CAXI4DMAIOI
<<
CAXI4DMAIlII
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
(
1
+
CAXI4DMAIOI
)
<<
CAXI4DMAIlII
)
)
)
begin
CAXI4DMAOl0I
=
CAXI4DMAIOI
;
end
else
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
127
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
128
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
127
;
end
else
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
63
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
64
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
63
;
end
else
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
31
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
32
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
31
;
end
else
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
15
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
16
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
15
;
end
else
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
7
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
8
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
7
;
end
else
if
(
(
CAXI4DMAIIOl
>=
(
1
+
(
3
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAlOOl
[
11
:
0
]
<=
13
'd
4096
-
(
4
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAOl0I
=
8
'd
3
;
end
else
begin
CAXI4DMAOl0I
=
8
'd
0
;
end
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAl0Il
==
1
'b
1
)
)
begin
CAXI4DMAl1II
=
1
'b
0
;
CAXI4DMAIOlI
=
32
'b
0
;
CAXI4DMAlIlI
=
2
'b
0
;
CAXI4DMAIllI
=
8
'b
0
;
CAXI4DMAOIlI
=
3
'b
0
;
CAXI4DMAl0II
=
CAXI4DMAOO1l
;
end
else
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAIOlI
=
CAXI4DMAlOOl
;
CAXI4DMAlIlI
=
CAXI4DMAlIOl
;
CAXI4DMAIllI
=
CAXI4DMAOl0I
;
CAXI4DMAOIlI
=
CAXI4DMAIlII
;
CAXI4DMAl0II
=
CAXI4DMAII0l
;
end
end
CAXI4DMAO00l
:
begin
if
(
CAXI4DMAll1
&
CAXI4DMAOll
)
begin
CAXI4DMAIOlI
=
32
'b
0
;
CAXI4DMAIllI
=
8
'b
0
;
CAXI4DMAOIlI
=
3
'b
0
;
CAXI4DMAlIlI
=
2
'b
0
;
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAl0Il
==
1
'b
1
)
)
begin
CAXI4DMAI1lI
=
{
{
(
AXI_DMA_DWIDTH
-
4
)
{
1
'b
0
}
}
,
1
'b
1
,
1
'b
0
,
CAXI4DMAOlI
[
1
:
0
]
}
;
CAXI4DMAlO0I
=
{
{
(
(
AXI_DMA_DWIDTH
/
8
)
-
1
)
{
1
'b
0
}
}
,
1
'b
1
}
;
end
else
begin
CAXI4DMAI1lI
=
{
{
(
AXI_DMA_DWIDTH
-
16
)
{
1
'b
0
}
}
,
CAXI4DMAO1I
,
{
8
{
1
'b
0
}
}
}
;
CAXI4DMAlO0I
=
{
{
(
(
AXI_DMA_DWIDTH
/
8
)
-
2
)
{
1
'b
0
}
}
,
1
'b
1
,
1
'b
0
}
;
end
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAOO0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAI00l
;
end
else
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAO00l
;
end
end
CAXI4DMAI00l
:
begin
if
(
CAXI4DMAO01
&
CAXI4DMAIll
)
begin
CAXI4DMAlO0I
=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
0
}
}
;
CAXI4DMAI1lI
=
{
AXI_DMA_DWIDTH
{
1
'b
0
}
}
;
CAXI4DMAOO0I
=
1
'b
0
;
CAXI4DMAII0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAl00l
;
end
else
begin
CAXI4DMAl0lI
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAI00l
;
end
end
CAXI4DMAl00l
:
begin
if
(
CAXI4DMAlll
&
CAXI4DMAl01
)
begin
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAl0Il
==
1
'b
1
)
)
begin
CAXI4DMAO1Il
=
1
'b
0
;
CAXI4DMAI00
=
1
'b
1
;
end
else
begin
CAXI4DMAO0Ol
=
1
'b
1
;
end
CAXI4DMAl0II
=
CAXI4DMAOI0l
;
end
else
begin
CAXI4DMAII0I
=
1
'b
1
;
CAXI4DMAl0II
=
CAXI4DMAl00l
;
end
end
CAXI4DMAOO1l
:
begin
if
(
CAXI4DMAOIOl
<
(
(
CAXI4DMAOllI
+
1
)
<<
CAXI4DMAIlII
)
)
begin
CAXI4DMAlOll
=
(
(
CAXI4DMAII1I
<<
CAXI4DMAIlII
)
+
(
CAXI4DMAOIOl
[
CAXI4DMAIlII
-
1
:
0
]
)
)
;
end
else
begin
CAXI4DMAlOll
=
(
(
CAXI4DMAOllI
+
1
)
<<
CAXI4DMAIlII
)
;
end
CAXI4DMAl0II
=
CAXI4DMAl10l
;
end
CAXI4DMAl10l
:
begin
if
(
CAXI4DMAIOl
>=
CAXI4DMAIOll
)
begin
CAXI4DMAl1II
=
1
'b
1
;
CAXI4DMAIOlI
=
CAXI4DMAIOOl
;
CAXI4DMAOIlI
=
CAXI4DMAIlII
;
CAXI4DMAIllI
=
CAXI4DMAlI0I
;
CAXI4DMAlIlI
=
CAXI4DMAlIOl
;
CAXI4DMAl0II
=
CAXI4DMAII0l
;
end
else
begin
CAXI4DMAl0II
=
CAXI4DMAl10l
;
end
end
default
:
begin
CAXI4DMAl0II
=
CAXI4DMAOI0l
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI0I
<=
8
'b
0
;
end
else
begin
CAXI4DMAlI0I
<=
CAXI4DMAOl0I
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlIOl
<=
2
'b
0
;
end
else
begin
CAXI4DMAlIOl
<=
CAXI4DMAOlOl
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIOOl
<=
32
'b
0
;
end
else
begin
CAXI4DMAIOOl
<=
CAXI4DMAlOOl
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIOl
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAOIOl
<=
CAXI4DMAIIOl
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1II
<=
1
'b
0
;
end
else
begin
CAXI4DMAI1II
<=
CAXI4DMAl1II
;
end
end
assign
CAXI4DMAll1
=
CAXI4DMAI1II
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOOlI
<=
32
'b
0
;
end
else
begin
CAXI4DMAOOlI
<=
CAXI4DMAIOlI
;
end
end
assign
CAXI4DMAl11
=
CAXI4DMAOOlI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlOlI
<=
3
'b
0
;
end
else
begin
CAXI4DMAlOlI
<=
CAXI4DMAOIlI
;
end
end
assign
CAXI4DMAlOOI
=
CAXI4DMAlOlI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIIlI
<=
2
'b
0
;
end
else
begin
CAXI4DMAIIlI
<=
CAXI4DMAlIlI
;
end
end
assign
CAXI4DMAOIOI
=
CAXI4DMAIIlI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOllI
<=
8
'b
0
;
end
else
begin
CAXI4DMAOllI
<=
CAXI4DMAIllI
;
end
end
assign
CAXI4DMAIOOI
=
CAXI4DMAOllI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlllI
<=
{
ID_WIDTH
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAlllI
<=
CAXI4DMAO0lI
;
end
end
assign
CAXI4DMAOOOI
=
CAXI4DMAlllI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI0lI
<=
1
'b
0
;
end
else
begin
CAXI4DMAI0lI
<=
CAXI4DMAl0lI
;
end
end
assign
CAXI4DMAO01
=
CAXI4DMAI0lI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO1lI
<=
{
AXI_DMA_DWIDTH
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAO1lI
<=
CAXI4DMAI1lI
;
end
end
assign
CAXI4DMAlIOI
=
CAXI4DMAO1lI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl1lI
<=
1
'b
0
;
end
else
begin
CAXI4DMAl1lI
<=
CAXI4DMAOO0I
;
end
end
assign
CAXI4DMAI01
=
CAXI4DMAl1lI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO0I
<=
{
(
AXI_DMA_DWIDTH
/
8
)
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIO0I
<=
CAXI4DMAlO0I
;
end
end
assign
CAXI4DMAIIOI
=
CAXI4DMAIO0I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOI0I
<=
1
'b
0
;
end
else
begin
CAXI4DMAOI0I
<=
CAXI4DMAII0I
;
end
end
assign
CAXI4DMAl01
=
CAXI4DMAOI0I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlIIl
<=
1
'b
0
;
end
else
begin
CAXI4DMAlIIl
<=
CAXI4DMAOlIl
;
end
end
assign
CAXI4DMAIO1l
=
CAXI4DMAlIIl
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIlIl
<=
{
CAXI4DMAOlII
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIlIl
<=
CAXI4DMAllIl
;
end
end
assign
CAXI4DMAOl1
=
CAXI4DMAIlIl
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO00I
<=
8
'b
0
;
end
else
begin
CAXI4DMAO00I
<=
CAXI4DMAI00I
;
end
end
assign
CAXI4DMAlI1
=
CAXI4DMAO00I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIl0I
<=
9
'b
0
;
end
else
begin
CAXI4DMAIl0I
<=
CAXI4DMAll0I
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIlOl
<=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIlOl
<=
CAXI4DMAllOl
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0Il
<=
1
'b
0
;
end
else
begin
CAXI4DMAl0Il
<=
CAXI4DMAO1Il
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl1Il
<=
1
'b
0
;
end
else
begin
CAXI4DMAl1Il
<=
CAXI4DMAOOll
;
end
end
assign
CAXI4DMAOl0
=
CAXI4DMAl1Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIOll
<=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIOll
<=
CAXI4DMAlOll
;
end
end
assign
CAXI4DMAIl0
=
CAXI4DMAIOll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAllII
<=
CAXI4DMAlIll
;
end
else
begin
CAXI4DMAllII
<=
CAXI4DMAO0II
;
end
end
always
@
(
*
)
begin
CAXI4DMAO10I
<=
1
'b
0
;
CAXI4DMAl10I
<=
CAXI4DMAI10I
;
CAXI4DMAl01I
<=
{
ID_WIDTH
{
1
'b
0
}
}
;
CAXI4DMAlI1I
<=
CAXI4DMAII1I
;
CAXI4DMAIO1I
<=
CAXI4DMAOO1I
;
CAXI4DMAOI1I
<=
CAXI4DMAlO1I
;
CAXI4DMAIl1I
<=
1
'b
0
;
CAXI4DMAOOIl
<=
1
'b
0
;
CAXI4DMAO01I
<=
CAXI4DMAll1I
;
CAXI4DMAIIIl
<=
{
CAXI4DMAOlII
{
1
'b
0
}
}
;
CAXI4DMAlOIl
<=
{
AXI_DMA_DWIDTH
{
1
'b
0
}
}
;
CAXI4DMAl1l
<=
1
'b
0
;
CAXI4DMAIO0
<=
1
'b
0
;
CAXI4DMAlI0
<=
{
CAXI4DMAO1OI
{
1
'b
0
}
}
;
CAXI4DMAII0
<=
1
'b
0
;
CAXI4DMAI11I
<=
CAXI4DMAO11I
;
CAXI4DMAOOOl
<=
CAXI4DMAl11I
;
CAXI4DMAI0Ol
<=
1
'b
0
;
CAXI4DMAl0Ol
<=
CAXI4DMAI10
;
CAXI4DMAO1Ol
<=
CAXI4DMAl10
;
CAXI4DMAI1Ol
<=
CAXI4DMAO10
;
CAXI4DMAI0Il
<=
CAXI4DMAO0Il
;
CAXI4DMAOIll
<=
1
'b
0
;
CAXI4DMAIIll
<=
1
'b
0
;
case
(
CAXI4DMAllII
)
CAXI4DMAlIll
:
begin
if
(
CAXI4DMAII
)
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAl10I
<=
CAXI4DMAIl
;
CAXI4DMAIO1I
<=
CAXI4DMAIlII
;
if
(
CAXI4DMAlI
==
2
'b
10
)
begin
CAXI4DMAOI1I
<=
2
'b
00
;
end
else
begin
CAXI4DMAOI1I
<=
2
'b
01
;
end
if
(
(
CAXI4DMAOl
>=
(
1
+
(
CAXI4DMAO0
<<
CAXI4DMAIlII
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
(
1
+
CAXI4DMAO0
)
<<
CAXI4DMAIlII
)
)
)
begin
CAXI4DMAlI1I
<=
CAXI4DMAO0
;
CAXI4DMAI11I
<=
CAXI4DMAO0
;
end
else
if
(
(
CAXI4DMAOl
>=
(
1
+
(
127
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
128
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAlI1I
<=
8
'd
127
;
CAXI4DMAI11I
<=
8
'd
127
;
end
else
if
(
(
CAXI4DMAOl
>=
(
1
+
(
63
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
64
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAlI1I
<=
8
'd
63
;
CAXI4DMAI11I
<=
8
'd
63
;
end
else
if
(
(
CAXI4DMAOl
>=
(
1
+
(
31
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
32
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAlI1I
<=
8
'd
31
;
CAXI4DMAI11I
<=
8
'd
31
;
end
else
if
(
(
CAXI4DMAOl
>=
(
1
+
(
15
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
16
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAlI1I
<=
8
'd
15
;
CAXI4DMAI11I
<=
8
'd
15
;
end
else
if
(
(
CAXI4DMAOl
>=
(
1
+
(
7
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
8
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAlI1I
<=
8
'd
7
;
CAXI4DMAI11I
<=
8
'd
7
;
end
else
if
(
(
CAXI4DMAOl
>=
(
1
+
(
3
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
&&
(
CAXI4DMAIl
[
11
:
0
]
<=
13
'd
4096
-
(
4
*
(
AXI_DMA_DWIDTH
/
8
)
)
)
)
begin
CAXI4DMAlI1I
<=
8
'd
3
;
CAXI4DMAI11I
<=
8
'd
3
;
end
else
begin
CAXI4DMAlI1I
<=
8
'd
0
;
CAXI4DMAI11I
<=
8
'd
0
;
end
CAXI4DMAOOOl
<=
CAXI4DMAOl
;
CAXI4DMAO0II
<=
CAXI4DMAOlll
;
end
else
if
(
CAXI4DMAllI
)
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAl10I
<=
CAXI4DMAI0I
;
CAXI4DMAIO1I
<=
CAXI4DMAIlII
;
CAXI4DMAOI1I
<=
2
'b
01
;
CAXI4DMAO0II
<=
CAXI4DMAI0ll
;
if
(
AXI_DMA_DWIDTH
==
32
)
begin
CAXI4DMAlI1I
<=
8
'd
4
;
end
else
if
(
AXI_DMA_DWIDTH
==
64
)
begin
CAXI4DMAlI1I
<=
8
'd
2
;
end
else
if
(
AXI_DMA_DWIDTH
==
128
)
begin
CAXI4DMAlI1I
<=
8
'd
1
;
end
else
begin
CAXI4DMAlI1I
<=
8
'd
0
;
end
end
else
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAIlI
)
)
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAl10I
<=
CAXI4DMAI0I
;
CAXI4DMAIO1I
<=
CAXI4DMAIlII
;
CAXI4DMAOI1I
<=
2
'b
01
;
CAXI4DMAO0II
<=
CAXI4DMAIO0l
;
if
(
AXI_DMA_DWIDTH
==
32
)
begin
CAXI4DMAlI1I
<=
8
'd
2
;
end
else
if
(
AXI_DMA_DWIDTH
==
64
)
begin
CAXI4DMAlI1I
<=
8
'd
1
;
end
else
begin
CAXI4DMAlI1I
<=
8
'd
0
;
end
end
else
if
(
CAXI4DMAO0I
)
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAl10I
<=
CAXI4DMAI0I
;
CAXI4DMAlI1I
<=
8
'd
0
;
CAXI4DMAIO1I
<=
CAXI4DMAIlII
;
CAXI4DMAOI1I
<=
2
'b
01
;
CAXI4DMAO0II
<=
CAXI4DMAO1ll
;
end
else
if
(
(
AXI4_STREAM_IF
==
1
)
&&
(
CAXI4DMAlOI
==
1
'b
1
)
)
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAl10I
<=
CAXI4DMAOII
;
CAXI4DMAlI1I
<=
8
'd
0
;
CAXI4DMAIO1I
<=
CAXI4DMAIlII
;
CAXI4DMAOI1I
<=
2
'b
01
;
CAXI4DMAO0II
<=
CAXI4DMAl1ll
;
end
else
begin
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
end
end
CAXI4DMAOlll
:
begin
if
(
CAXI4DMAO11
&
CAXI4DMAO0l
)
begin
CAXI4DMAl10I
<=
32
'b
0
;
CAXI4DMAlI1I
<=
8
'b
0
;
CAXI4DMAIO1I
<=
3
'b
0
;
CAXI4DMAOI1I
<=
2
'b
0
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAIlll
;
if
(
CAXI4DMAl11I
<
(
(
CAXI4DMAII1I
+
1
)
<<
CAXI4DMAIlII
)
)
begin
CAXI4DMAlI0
<=
(
(
CAXI4DMAII1I
<<
CAXI4DMAIlII
)
+
(
CAXI4DMAl11I
[
CAXI4DMAIlII
-
1
:
0
]
)
)
;
end
else
begin
CAXI4DMAlI0
<=
(
(
CAXI4DMAII1I
+
1
)
<<
CAXI4DMAIlII
)
;
end
CAXI4DMAII0
<=
1
'b
1
;
end
else
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAOlll
;
end
end
CAXI4DMAIlll
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
)
begin
CAXI4DMAOOIl
<=
1
'b
1
;
CAXI4DMAlOIl
<=
CAXI4DMAIIl
;
if
(
CAXI4DMAO1l
)
begin
if
(
CAXI4DMAl11I
<
(
(
CAXI4DMAO11I
+
1
)
<<
CAXI4DMAIlII
)
)
begin
CAXI4DMAIIIl
<=
{
1
'b
0
,
CAXI4DMAl11I
[
CAXI4DMAIlII
-
1
:
0
]
}
;
end
else
begin
CAXI4DMAIIIl
<=
(
AXI_DMA_DWIDTH
/
8
)
;
end
CAXI4DMAO0II
<=
CAXI4DMAO0ll
;
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAIIIl
<=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAO0II
<=
CAXI4DMAllll
;
end
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAIlll
;
end
end
CAXI4DMAllll
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
)
begin
CAXI4DMAOOIl
<=
1
'b
1
;
CAXI4DMAlOIl
<=
CAXI4DMAIIl
;
CAXI4DMAO01I
<=
CAXI4DMAll1I
+
1
'b
1
;
if
(
CAXI4DMAO1l
)
begin
if
(
CAXI4DMAl11I
<
(
(
CAXI4DMAO11I
+
1
)
<<
CAXI4DMAIlII
)
)
begin
CAXI4DMAIIIl
<=
{
1
'b
0
,
CAXI4DMAl11I
[
CAXI4DMAIlII
-
1
:
0
]
}
;
end
else
begin
CAXI4DMAIIIl
<=
(
AXI_DMA_DWIDTH
/
8
)
;
end
CAXI4DMAO0II
<=
CAXI4DMAO0ll
;
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAIIIl
<=
(
AXI_DMA_DWIDTH
/
8
)
;
CAXI4DMAO0II
<=
CAXI4DMAllll
;
end
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAllll
;
end
end
CAXI4DMAO0ll
:
begin
CAXI4DMAO01I
<=
8
'b
0
;
CAXI4DMAl1l
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
end
CAXI4DMAI0ll
:
begin
if
(
CAXI4DMAO11
&
CAXI4DMAO0l
)
begin
CAXI4DMAl10I
<=
32
'b
0
;
CAXI4DMAlI1I
<=
8
'b
0
;
CAXI4DMAIO1I
<=
3
'b
0
;
CAXI4DMAOI1I
<=
2
'b
0
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAl0ll
;
end
else
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAI0ll
;
end
end
CAXI4DMAl0ll
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
)
begin
if
(
CAXI4DMAO1l
)
begin
CAXI4DMAI0Il
<=
2
'b
0
;
CAXI4DMAI0Ol
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
if
(
(
AXI_DMA_DWIDTH
==
256
)
||
(
AXI_DMA_DWIDTH
==
512
)
)
begin
CAXI4DMAl0Ol
[
133
:
0
]
<=
{
CAXI4DMAIIl
[
159
:
64
]
,
CAXI4DMAIIl
[
55
:
32
]
,
CAXI4DMAIIl
[
13
:
0
]
}
;
CAXI4DMAI1Ol
<=
{
CAXI4DMAIIl
[
14
]
,
CAXI4DMAIIl
[
13
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
15
]
;
end
else
begin
CAXI4DMAl0Ol
[
133
:
102
]
<=
CAXI4DMAIIl
[
31
:
0
]
;
CAXI4DMAl0Ol
[
101
:
0
]
<=
CAXI4DMAI10
[
101
:
0
]
;
end
end
else
begin
CAXI4DMAI0Il
<=
CAXI4DMAO0Il
+
1
'b
1
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAl0ll
;
if
(
AXI_DMA_DWIDTH
==
64
)
begin
if
(
CAXI4DMAO0Il
==
2
'd
1
)
begin
CAXI4DMAl0Ol
[
133
:
102
]
<=
CAXI4DMAI10
[
133
:
102
]
;
CAXI4DMAl0Ol
[
101
:
38
]
<=
CAXI4DMAIIl
[
63
:
0
]
;
CAXI4DMAl0Ol
[
37
:
0
]
<=
CAXI4DMAI10
[
37
:
0
]
;
end
else
begin
CAXI4DMAl0Ol
[
133
:
38
]
<=
CAXI4DMAI10
[
133
:
38
]
;
CAXI4DMAl0Ol
[
37
:
0
]
<=
{
CAXI4DMAIIl
[
55
:
32
]
,
CAXI4DMAIIl
[
13
:
0
]
}
;
CAXI4DMAI1Ol
<=
{
CAXI4DMAIIl
[
14
]
,
CAXI4DMAIIl
[
13
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
15
]
;
end
end
else
if
(
AXI_DMA_DWIDTH
==
128
)
begin
CAXI4DMAl0Ol
[
133
:
102
]
<=
CAXI4DMAI10
[
133
:
102
]
;
CAXI4DMAl0Ol
[
101
:
0
]
<=
{
CAXI4DMAIIl
[
127
:
64
]
,
CAXI4DMAIIl
[
55
:
32
]
,
CAXI4DMAIIl
[
13
:
0
]
}
;
CAXI4DMAI1Ol
<=
{
CAXI4DMAIIl
[
14
]
,
CAXI4DMAIIl
[
13
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
15
]
;
end
else
begin
if
(
CAXI4DMAO0Il
==
2
'd
1
)
begin
CAXI4DMAl0Ol
[
133
:
38
]
<=
CAXI4DMAI10
[
133
:
38
]
;
CAXI4DMAl0Ol
[
37
:
14
]
<=
CAXI4DMAIIl
[
23
:
0
]
;
CAXI4DMAl0Ol
[
13
:
0
]
<=
CAXI4DMAI10
[
13
:
0
]
;
end
else
if
(
CAXI4DMAO0Il
==
2
'd
2
)
begin
CAXI4DMAl0Ol
[
133
:
70
]
<=
CAXI4DMAI10
[
133
:
70
]
;
CAXI4DMAl0Ol
[
69
:
38
]
<=
CAXI4DMAIIl
[
31
:
0
]
;
CAXI4DMAl0Ol
[
37
:
0
]
<=
CAXI4DMAI10
[
37
:
0
]
;
end
else
if
(
CAXI4DMAO0Il
==
2
'd
3
)
begin
CAXI4DMAl0Ol
[
133
:
102
]
<=
CAXI4DMAI10
[
133
:
102
]
;
CAXI4DMAl0Ol
[
101
:
70
]
<=
CAXI4DMAIIl
[
31
:
0
]
;
CAXI4DMAl0Ol
[
69
:
0
]
<=
CAXI4DMAI10
[
69
:
0
]
;
end
else
begin
CAXI4DMAl0Ol
[
133
:
14
]
<=
CAXI4DMAI10
[
133
:
14
]
;
CAXI4DMAl0Ol
[
13
:
0
]
<=
CAXI4DMAIIl
[
13
:
0
]
;
CAXI4DMAI1Ol
<=
{
CAXI4DMAIIl
[
14
]
,
CAXI4DMAIIl
[
13
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
15
]
;
end
end
end
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAl0ll
;
end
end
CAXI4DMAO1ll
:
begin
if
(
CAXI4DMAO11
&
CAXI4DMAO0l
)
begin
CAXI4DMAl10I
<=
32
'b
0
;
CAXI4DMAlI1I
<=
8
'b
0
;
CAXI4DMAIO1I
<=
3
'b
0
;
CAXI4DMAOI1I
<=
2
'b
0
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAI1ll
;
end
else
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAO1ll
;
end
end
CAXI4DMAI1ll
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
&
CAXI4DMAO1l
)
begin
CAXI4DMAI0Ol
<=
1
'b
1
;
CAXI4DMAI1Ol
<=
{
CAXI4DMAIIl
[
14
]
,
CAXI4DMAIIl
[
13
]
}
;
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAI1ll
;
end
end
CAXI4DMAl1ll
:
begin
if
(
CAXI4DMAO11
&
CAXI4DMAO0l
)
begin
CAXI4DMAl10I
<=
32
'b
0
;
CAXI4DMAlI1I
<=
8
'b
0
;
CAXI4DMAIO1I
<=
3
'b
0
;
CAXI4DMAOI1I
<=
2
'b
0
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAOO0l
;
end
else
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAl1ll
;
end
end
CAXI4DMAOO0l
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
&
CAXI4DMAO1l
)
begin
CAXI4DMAIIll
<=
CAXI4DMAIIl
[
2
]
;
CAXI4DMAOIll
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAOO0l
;
end
end
CAXI4DMAIO0l
:
begin
if
(
CAXI4DMAO11
&
CAXI4DMAO0l
)
begin
CAXI4DMAl10I
<=
32
'b
0
;
CAXI4DMAlI1I
<=
8
'b
0
;
CAXI4DMAIO1I
<=
3
'b
0
;
CAXI4DMAOI1I
<=
2
'b
0
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlO0l
;
end
else
begin
CAXI4DMAO10I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAIO0l
;
end
end
CAXI4DMAlO0l
:
begin
if
(
CAXI4DMAI0l
&
CAXI4DMAI11
)
begin
if
(
CAXI4DMAO1l
)
begin
CAXI4DMAI0Il
<=
2
'b
0
;
CAXI4DMAI0Ol
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
if
(
(
AXI_DMA_DWIDTH
==
128
)
||
(
AXI_DMA_DWIDTH
==
256
)
||
(
AXI_DMA_DWIDTH
==
512
)
)
begin
CAXI4DMAl0Ol
[
133
:
58
]
<=
{
76
{
1
'b
0
}
}
;
CAXI4DMAl0Ol
[
57
:
26
]
<=
CAXI4DMAIIl
[
95
:
64
]
;
CAXI4DMAl0Ol
[
25
:
2
]
<=
CAXI4DMAIIl
[
55
:
32
]
;
CAXI4DMAl0Ol
[
1
:
0
]
<=
CAXI4DMAIIl
[
1
:
0
]
;
CAXI4DMAI1Ol
<=
{
1
'b
0
,
CAXI4DMAIIl
[
2
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
3
]
;
end
else
begin
CAXI4DMAl0Ol
[
133
:
58
]
<=
{
76
{
1
'b
0
}
}
;
CAXI4DMAl0Ol
[
57
:
26
]
<=
CAXI4DMAIIl
[
31
:
0
]
;
CAXI4DMAl0Ol
[
25
:
0
]
<=
CAXI4DMAI10
[
25
:
0
]
;
end
end
else
begin
CAXI4DMAI0Il
<=
CAXI4DMAO0Il
+
1
'b
1
;
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlO0l
;
if
(
AXI_DMA_DWIDTH
==
64
)
begin
CAXI4DMAl0Ol
[
133
:
26
]
<=
{
108
{
1
'b
0
}
}
;
CAXI4DMAl0Ol
[
25
:
0
]
<=
{
CAXI4DMAIIl
[
55
:
32
]
,
CAXI4DMAIIl
[
1
:
0
]
}
;
CAXI4DMAI1Ol
<=
{
1
'b
0
,
CAXI4DMAIIl
[
2
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
3
]
;
end
else
begin
if
(
CAXI4DMAO0Il
==
2
'd
1
)
begin
CAXI4DMAl0Ol
[
133
:
26
]
<=
CAXI4DMAI10
[
133
:
26
]
;
CAXI4DMAl0Ol
[
25
:
2
]
<=
CAXI4DMAIIl
[
23
:
0
]
;
CAXI4DMAl0Ol
[
1
:
0
]
<=
CAXI4DMAI10
[
1
:
0
]
;
end
else
begin
CAXI4DMAl0Ol
[
133
:
2
]
<=
{
132
{
1
'b
0
}
}
;
CAXI4DMAl0Ol
[
1
:
0
]
<=
CAXI4DMAIIl
[
1
:
0
]
;
CAXI4DMAI1Ol
<=
{
1
'b
0
,
CAXI4DMAIIl
[
2
]
}
;
CAXI4DMAO1Ol
<=
CAXI4DMAIIl
[
3
]
;
end
end
end
end
else
begin
CAXI4DMAIl1I
<=
1
'b
1
;
CAXI4DMAO0II
<=
CAXI4DMAlO0l
;
end
end
default
:
begin
CAXI4DMAO0II
<=
CAXI4DMAlIll
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl11I
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAl11I
<=
CAXI4DMAOOOl
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO11I
<=
8
'b
0
;
end
else
begin
CAXI4DMAO11I
<=
CAXI4DMAI11I
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl00I
<=
1
'b
0
;
end
else
begin
CAXI4DMAl00I
<=
CAXI4DMAO10I
;
end
end
assign
CAXI4DMAO11
=
CAXI4DMAl00I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI10I
<=
32
'b
0
;
end
else
begin
CAXI4DMAI10I
<=
CAXI4DMAl10I
;
end
end
assign
CAXI4DMAOlOI
=
CAXI4DMAI10I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOO1I
<=
3
'b
0
;
end
else
begin
CAXI4DMAOO1I
<=
CAXI4DMAIO1I
;
end
end
assign
CAXI4DMAO0OI
=
CAXI4DMAOO1I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlO1I
<=
2
'b
0
;
end
else
begin
CAXI4DMAlO1I
<=
CAXI4DMAOI1I
;
end
end
assign
CAXI4DMAI0OI
=
CAXI4DMAlO1I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI01I
<=
{
ID_WIDTH
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAI01I
<=
CAXI4DMAl01I
;
end
end
assign
CAXI4DMAIlOI
=
CAXI4DMAI01I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAII1I
<=
8
'b
0
;
end
else
begin
CAXI4DMAII1I
<=
CAXI4DMAlI1I
;
end
end
assign
CAXI4DMAllOI
=
CAXI4DMAII1I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOl1I
<=
1
'b
0
;
end
else
begin
CAXI4DMAOl1I
<=
CAXI4DMAIl1I
;
end
end
assign
CAXI4DMAI11
=
CAXI4DMAOl1I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAll1I
<=
8
'b
0
;
end
else
begin
CAXI4DMAll1I
<=
CAXI4DMAO01I
;
end
end
assign
CAXI4DMAIO1
=
CAXI4DMAll1I
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI10
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAI10
<=
CAXI4DMAl0Ol
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10
<=
1
'b
0
;
end
else
begin
CAXI4DMAl10
<=
CAXI4DMAO1Ol
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl00
<=
1
'b
0
;
end
else
begin
CAXI4DMAl00
<=
CAXI4DMAO0Ol
|
CAXI4DMAI0Ol
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO10
<=
2
'b
0
;
end
else
begin
CAXI4DMAO10
<=
CAXI4DMAI1Ol
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl1Ol
<=
1
'b
0
;
end
else
begin
CAXI4DMAl1Ol
<=
CAXI4DMAOOIl
;
end
end
assign
CAXI4DMAOO1
=
CAXI4DMAl1Ol
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIOIl
<=
{
AXI_DMA_DWIDTH
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIOIl
<=
CAXI4DMAlOIl
;
end
end
assign
CAXI4DMAlO1
=
CAXI4DMAIOIl
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIIl
<=
{
CAXI4DMAOlII
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAOIIl
<=
CAXI4DMAIIIl
;
end
end
assign
CAXI4DMAOI1
=
CAXI4DMAOIIl
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO0Il
<=
2
'b
0
;
end
else
begin
CAXI4DMAO0Il
<=
CAXI4DMAI0Il
;
end
end
assign
CAXI4DMAOI1
=
CAXI4DMAOIIl
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAll0
<=
1
'b
0
;
end
else
begin
CAXI4DMAll0
<=
CAXI4DMAOIll
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO00
<=
1
'b
0
;
end
else
begin
CAXI4DMAO00
<=
CAXI4DMAIIll
;
end
end
endmodule
