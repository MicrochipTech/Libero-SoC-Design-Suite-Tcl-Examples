// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAO0I1I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAIll0I
,
CAXI4DMAl0l0I
,
CAXI4DMAl0I1I
,
CAXI4DMAO0l0I
,
CAXI4DMAO1l0I
,
CAXI4DMAOO10I
,
CAXI4DMAIO10I
,
CAXI4DMAlO10I
,
CAXI4DMAOI10I
,
CAXI4DMAO1I0I
,
CAXI4DMAO1I1I
,
CAXI4DMAI1O1I
,
CAXI4DMAOIllI
,
valid
,
CAXI4DMAlIlOI
,
CAXI4DMAOllOI
,
CAXI4DMAIllOI
,
CAXI4DMAlllOI
,
intDscrptrNum
,
CAXI4DMAII0OI
,
CAXI4DMAlI0OI
,
strDscrptr
,
CAXI4DMAI1I1I
,
CAXI4DMAI1I0I
)
;
parameter
CAXI4DMAOIO1
=
2
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAIll0I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl0l0I
;
input
CAXI4DMAl0I1I
;
input
CAXI4DMAO0l0I
;
input
[
31
:
0
]
CAXI4DMAO1l0I
;
input
CAXI4DMAOO10I
;
input
CAXI4DMAIO10I
;
input
CAXI4DMAlO10I
;
input
CAXI4DMAOI10I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO1I0I
;
input
CAXI4DMAO1I1I
;
input
[
31
:
0
]
CAXI4DMAI1O1I
;
input
CAXI4DMAOIllI
;
output
reg
valid
;
output
reg
CAXI4DMAlIlOI
;
output
reg
CAXI4DMAOllOI
;
output
reg
CAXI4DMAIllOI
;
output
reg
CAXI4DMAlllOI
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
intDscrptrNum
;
output
reg
CAXI4DMAII0OI
;
output
reg
[
31
:
0
]
CAXI4DMAlI0OI
;
output
reg
strDscrptr
;
output
reg
CAXI4DMAI1I1I
;
output
reg
CAXI4DMAI1I0I
;
reg
[
1
:
0
]
CAXI4DMAl10OI
;
reg
[
1
:
0
]
CAXI4DMAOO1OI
;
localparam
[
1
:
0
]
CAXI4DMAO0O0l
=
2
'b
01
;
localparam
[
1
:
0
]
CAXI4DMAI0O0l
=
2
'b
10
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO0O0l
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
valid
<=
1
'b
0
;
CAXI4DMAlllOI
<=
1
'b
0
;
intDscrptrNum
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAlI0OI
<=
32
'b
0
;
CAXI4DMAI1I0I
<=
1
'b
0
;
CAXI4DMAlIlOI
<=
1
'b
0
;
CAXI4DMAOllOI
<=
1
'b
0
;
CAXI4DMAIllOI
<=
1
'b
0
;
CAXI4DMAI1I1I
<=
1
'b
0
;
CAXI4DMAII0OI
<=
1
'b
0
;
strDscrptr
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO0O0l
:
begin
if
(
CAXI4DMAIll0I
)
begin
valid
<=
1
'b
1
;
CAXI4DMAlllOI
<=
1
'b
1
;
intDscrptrNum
<=
CAXI4DMAl0l0I
;
CAXI4DMAII0OI
<=
CAXI4DMAl0I1I
;
strDscrptr
<=
CAXI4DMAO0l0I
;
CAXI4DMAlI0OI
<=
CAXI4DMAO1l0I
;
CAXI4DMAI1I0I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI0O0l
;
end
else
if
(
CAXI4DMAOO10I
)
begin
valid
<=
1
'b
1
;
CAXI4DMAlIlOI
<=
CAXI4DMAIO10I
;
CAXI4DMAOllOI
<=
CAXI4DMAlO10I
;
CAXI4DMAIllOI
<=
CAXI4DMAOI10I
;
intDscrptrNum
<=
CAXI4DMAO1I0I
;
CAXI4DMAII0OI
<=
CAXI4DMAO1I1I
;
CAXI4DMAlI0OI
<=
CAXI4DMAI1O1I
;
strDscrptr
<=
CAXI4DMAOIllI
;
CAXI4DMAI1I1I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO0O0l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO0O0l
;
end
end
CAXI4DMAI0O0l
:
begin
if
(
CAXI4DMAOO10I
)
begin
valid
<=
1
'b
1
;
CAXI4DMAlIlOI
<=
CAXI4DMAIO10I
;
CAXI4DMAOllOI
<=
CAXI4DMAlO10I
;
CAXI4DMAIllOI
<=
CAXI4DMAOI10I
;
intDscrptrNum
<=
CAXI4DMAO1I0I
;
CAXI4DMAII0OI
<=
CAXI4DMAO1I1I
;
CAXI4DMAlI0OI
<=
CAXI4DMAI1O1I
;
strDscrptr
<=
CAXI4DMAOIllI
;
CAXI4DMAI1I1I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO0O0l
;
end
else
if
(
CAXI4DMAIll0I
)
begin
valid
<=
1
'b
1
;
CAXI4DMAlllOI
<=
1
'b
1
;
intDscrptrNum
<=
CAXI4DMAl0l0I
;
strDscrptr
<=
CAXI4DMAO0l0I
;
CAXI4DMAII0OI
<=
CAXI4DMAl0I1I
;
CAXI4DMAlI0OI
<=
CAXI4DMAO1l0I
;
CAXI4DMAI1I0I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAI0O0l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAI0O0l
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO0O0l
;
end
endcase
end
endmodule
