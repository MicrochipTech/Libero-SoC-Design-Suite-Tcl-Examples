//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Sep  9 11:10:12 2020
// Version: v12.4 12.900.0.16
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// TOP
module TOP(
    // Inputs
    A,
    CLK,
    D,
    // Outputs
    Q
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  A;
input  CLK;
input  D;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Q;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   A;
wire   AND2_0_Y;
wire   CLK;
wire   D;
wire   DFN1_0_Q;
wire   Q_net_0;
wire   Q_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Q_net_1 = Q_net_0;
assign Q       = Q_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AND2
AND2 AND2_0(
        // Inputs
        .A ( A ),
        .B ( DFN1_0_Q ),
        // Outputs
        .Y ( AND2_0_Y ) 
        );

//--------DFN1
DFN1 DFN1_0(
        // Inputs
        .D   ( D ),
        .CLK ( CLK ),
        // Outputs
        .Q   ( DFN1_0_Q ) 
        );

//--------DFN1
DFN1 DFN1_1(
        // Inputs
        .D   ( AND2_0_Y ),
        .CLK ( CLK ),
        // Outputs
        .Q   ( Q_net_0 ) 
        );


endmodule
