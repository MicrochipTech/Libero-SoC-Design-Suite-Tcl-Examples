// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAII10
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAOO1
,
CAXI4DMAlO1
,
CAXI4DMAIO1l
,
CAXI4DMAI1Il
,
CAXI4DMAlI10
,
CAXI4DMAOl10
,
CAXI4DMAIl10
)
;
parameter
CAXI4DMAll10
=
8
;
parameter
CAXI4DMAO010
=
2
;
function
integer
CAXI4DMAIOII
;
input
integer
CAXI4DMAlOII
;
integer
CAXI4DMAOIII
,
CAXI4DMAIIII
,
CAXI4DMAlIII
;
begin
CAXI4DMAIIII
=
1
;
CAXI4DMAlIII
=
0
;
CAXI4DMAOIII
=
CAXI4DMAlOII
+
1
;
while
(
CAXI4DMAIIII
<
CAXI4DMAOIII
)
begin
CAXI4DMAIIII
=
CAXI4DMAIIII
*
2
;
CAXI4DMAlIII
=
CAXI4DMAlIII
+
1
;
end
CAXI4DMAIOII
=
CAXI4DMAlIII
;
end
endfunction
localparam
CAXI4DMAI010
=
CAXI4DMAO010
+
3
;
localparam
CAXI4DMAl010
=
CAXI4DMAIOII
(
CAXI4DMAI010
-
1
)
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAOO1
;
input
[
CAXI4DMAll10
-
1
:
0
]
CAXI4DMAlO1
;
input
CAXI4DMAIO1l
;
output
[
CAXI4DMAll10
-
1
:
0
]
CAXI4DMAI1Il
;
output
CAXI4DMAlI10
;
output
CAXI4DMAOl10
;
output
CAXI4DMAIl10
;
reg
[
CAXI4DMAll10
-
1
:
0
]
CAXI4DMAO110
[
0
:
CAXI4DMAI010
-
1
]
;
reg
[
CAXI4DMAl010
-
1
:
0
]
CAXI4DMAIO1
;
reg
[
CAXI4DMAl010
-
1
:
0
]
CAXI4DMAlI1
;
reg
[
CAXI4DMAl010
:
0
]
CAXI4DMAI110
;
always
@
(
posedge
CAXI4DMAI
)
begin
if
(
CAXI4DMAOO1
)
CAXI4DMAO110
[
CAXI4DMAIO1
]
<=
CAXI4DMAlO1
;
end
assign
CAXI4DMAI1Il
=
CAXI4DMAO110
[
CAXI4DMAlI1
]
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI110
<=
{
(
CAXI4DMAl010
+
1
)
{
1
'b
0
}
}
;
end
else
begin
case
(
{
CAXI4DMAOO1
,
CAXI4DMAIO1l
}
)
2
'b
01
:
begin
CAXI4DMAI110
<=
CAXI4DMAI110
-
1
'b
1
;
end
2
'b
10
:
begin
if
(
!
CAXI4DMAlI10
)
begin
CAXI4DMAI110
<=
CAXI4DMAI110
+
1
'b
1
;
end
else
begin
CAXI4DMAI110
<=
CAXI4DMAI110
;
end
end
default
:
begin
CAXI4DMAI110
<=
CAXI4DMAI110
;
end
endcase
end
end
assign
CAXI4DMAlI10
=
(
CAXI4DMAI110
==
CAXI4DMAI010
)
;
assign
CAXI4DMAIl10
=
(
CAXI4DMAI110
==
{
(
CAXI4DMAl010
+
1
)
{
1
'b
0
}
}
)
;
assign
CAXI4DMAOl10
=
(
CAXI4DMAI110
==
CAXI4DMAO010
)
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO1
<=
{
CAXI4DMAl010
{
1
'b
0
}
}
;
end
else
begin
if
(
CAXI4DMAOO1
)
begin
if
(
!
CAXI4DMAlI10
)
begin
CAXI4DMAIO1
<=
CAXI4DMAIO1
+
1
'b
1
;
end
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI1
<=
{
CAXI4DMAl010
{
1
'b
0
}
}
;
end
else
begin
if
(
CAXI4DMAIO1l
)
begin
CAXI4DMAlI1
<=
CAXI4DMAlI1
+
1
'b
1
;
end
end
end
endmodule
