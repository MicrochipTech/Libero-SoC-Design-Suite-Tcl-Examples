// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAl0IIl
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAOOOIl
,
CAXI4DMAlIOIl
,
strDscrptr
,
CAXI4DMAI1IlI
,
CAXI4DMAllllI
,
CAXI4DMAlOOIl
,
CAXI4DMAIIIIl
,
CAXI4DMAOIOIl
,
CAXI4DMAI1IIl
,
CAXI4DMAlI0OI
,
CAXI4DMAOO0Ol
,
CAXI4DMAl1IIl
,
CAXI4DMAOOlIl
,
CAXI4DMAIOlIl
,
CAXI4DMAlOlIl
,
CAXI4DMAOIlIl
,
CAXI4DMAIIlIl
,
CAXI4DMAlIlIl
,
CAXI4DMAOllIl
,
CAXI4DMAIllIl
,
CAXI4DMAlllIl
,
CAXI4DMAO0lIl
,
CAXI4DMAOO1Ol
,
CAXI4DMAI0lIl
,
CAXI4DMAOllOI
,
CAXI4DMAl0lIl
,
CAXI4DMAO1lIl
,
CAXI4DMAI10Ol
,
CAXI4DMAIOI
,
CAXI4DMAI0
,
CAXI4DMAlI0
,
CAXI4DMAOI
,
CAXI4DMAl0
,
CAXI4DMAI1
,
CAXI4DMAI101I
,
CAXI4DMAll
,
CAXI4DMAlOI
,
CAXI4DMAOII
,
CAXI4DMAl00Ol
)
;
parameter
NUM_PRI_LVLS
=
1
;
parameter
CAXI4DMAl0OI
=
0
;
parameter
CAXI4DMAO1OI
=
13
;
parameter
CAXI4DMAI1OI
=
8
;
parameter
PRI_0_NUM_OF_BEATS
=
255
;
parameter
PRI_1_NUM_OF_BEATS
=
127
;
parameter
PRI_2_NUM_OF_BEATS
=
63
;
parameter
PRI_3_NUM_OF_BEATS
=
31
;
parameter
PRI_4_NUM_OF_BEATS
=
15
;
parameter
PRI_5_NUM_OF_BEATS
=
7
;
parameter
PRI_6_NUM_OF_BEATS
=
3
;
parameter
PRI_7_NUM_OF_BEATS
=
0
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAOOOIl
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAlIOIl
;
input
strDscrptr
;
input
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAllllI
;
input
CAXI4DMAI1IlI
;
input
[
2
:
0
]
CAXI4DMAlOOIl
;
input
[
1
:
0
]
CAXI4DMAIIIIl
;
input
[
2
:
0
]
CAXI4DMAOIOIl
;
input
[
31
:
0
]
CAXI4DMAI1IIl
;
input
[
31
:
0
]
CAXI4DMAlI0OI
;
input
CAXI4DMAOO0Ol
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAl1IIl
;
input
CAXI4DMAOOlIl
;
input
CAXI4DMAIOlIl
;
input
CAXI4DMAlOlIl
;
input
CAXI4DMAOIlIl
;
input
CAXI4DMAIIlIl
;
input
CAXI4DMAlIlIl
;
input
CAXI4DMAOllIl
;
input
CAXI4DMAIllIl
;
input
CAXI4DMAlllIl
;
input
CAXI4DMAO0lIl
;
input
CAXI4DMAOO1Ol
;
output
CAXI4DMAI0lIl
;
output
CAXI4DMAOllOI
;
output
CAXI4DMAl0lIl
;
output
CAXI4DMAO1lIl
;
output
CAXI4DMAI10Ol
;
output
CAXI4DMAOI
;
output
[
1
:
0
]
CAXI4DMAl0
;
output
[
2
:
0
]
CAXI4DMAI1
;
output
[
31
:
0
]
CAXI4DMAI101I
;
output
[
2
:
0
]
CAXI4DMAll
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAlI0
;
output
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAIOI
;
output
CAXI4DMAI0
;
output
reg
CAXI4DMAlOI
;
output
reg
[
31
:
0
]
CAXI4DMAOII
;
output
CAXI4DMAl00Ol
;
reg
[
8
:
0
]
CAXI4DMAl10OI
;
reg
[
8
:
0
]
CAXI4DMAOO1OI
;
reg
CAXI4DMAIll1l
;
reg
CAXI4DMAlll1l
;
reg
CAXI4DMAlO0ll
;
reg
CAXI4DMAOI0ll
;
reg
CAXI4DMAO0l1l
;
reg
CAXI4DMAI0l1l
;
reg
CAXI4DMAl0l1l
;
reg
CAXI4DMAO1l1l
;
reg
CAXI4DMAI1l1l
;
reg
CAXI4DMAl1l1l
;
reg
[
31
:
0
]
CAXI4DMAOO01l
;
reg
[
31
:
0
]
CAXI4DMAIO01l
;
reg
[
1
:
0
]
CAXI4DMAlO01l
;
reg
[
1
:
0
]
CAXI4DMAOI01l
;
reg
[
2
:
0
]
CAXI4DMAII01l
;
reg
[
2
:
0
]
CAXI4DMAlI01l
;
reg
[
2
:
0
]
CAXI4DMAO1l0l
;
reg
[
2
:
0
]
CAXI4DMAI1l0l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAlI0Ol
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOl01l
;
reg
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAIl01l
;
reg
[
CAXI4DMAI1OI
-
1
:
0
]
CAXI4DMAll01l
;
reg
CAXI4DMAl0Il
;
reg
CAXI4DMAO1Il
;
reg
CAXI4DMAO001l
;
reg
CAXI4DMAI001l
;
reg
CAXI4DMAl001l
;
reg
CAXI4DMAO101l
;
localparam
[
8
:
0
]
CAXI4DMAO1OII
=
9
'b
000000001
;
localparam
[
8
:
0
]
CAXI4DMAI101l
=
9
'b
000000010
;
localparam
[
8
:
0
]
CAXI4DMAI000l
=
9
'b
000000100
;
localparam
[
8
:
0
]
CAXI4DMAl101l
=
9
'b
000001000
;
localparam
[
8
:
0
]
CAXI4DMAOO11l
=
9
'b
000010000
;
localparam
[
8
:
0
]
CAXI4DMAIO11l
=
9
'b
000100000
;
localparam
[
8
:
0
]
CAXI4DMAlO11l
=
9
'b
001000000
;
localparam
[
8
:
0
]
CAXI4DMAOI11l
=
9
'b
010000000
;
localparam
[
8
:
0
]
CAXI4DMAOO10l
=
9
'b
100000000
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAl1l1l
<=
1
'b
0
;
CAXI4DMAIO01l
<=
32
'b
0
;
CAXI4DMAOI01l
<=
2
'b
0
;
CAXI4DMAlI01l
<=
3
'b
0
;
CAXI4DMAI1l0l
<=
3
'b
0
;
CAXI4DMAlll1l
<=
1
'b
0
;
CAXI4DMAOI0ll
<=
1
'b
0
;
CAXI4DMAI0l1l
<=
1
'b
0
;
CAXI4DMAO1l1l
<=
1
'b
0
;
CAXI4DMAOl01l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAll01l
<=
CAXI4DMAIl01l
;
CAXI4DMAO1Il
<=
1
'b
0
;
CAXI4DMAlOI
<=
1
'b
0
;
CAXI4DMAOII
<=
32
'b
0
;
CAXI4DMAI001l
<=
1
'b
0
;
CAXI4DMAO101l
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAOOOIl
)
begin
if
(
CAXI4DMAIIIIl
==
2
'b
00
)
begin
CAXI4DMAO101l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO10l
;
end
else
if
(
strDscrptr
)
begin
if
(
CAXI4DMAI1IlI
==
1
'b
1
)
begin
CAXI4DMAl1l1l
<=
1
'b
1
;
CAXI4DMAO1Il
<=
1
'b
1
;
CAXI4DMAOl01l
<=
CAXI4DMAlIOIl
;
CAXI4DMAIO01l
<=
CAXI4DMAI1IIl
;
CAXI4DMAOI01l
<=
CAXI4DMAIIIIl
;
CAXI4DMAll01l
<=
PRI_0_NUM_OF_BEATS
;
CAXI4DMAOO1OI
<=
CAXI4DMAI101l
;
end
else
begin
CAXI4DMAlOI
<=
1
'b
1
;
CAXI4DMAOII
<=
CAXI4DMAlI0OI
;
CAXI4DMAOO1OI
<=
CAXI4DMAOI11l
;
end
end
else
if
(
CAXI4DMAOO0Ol
)
begin
CAXI4DMAl1l1l
<=
1
'b
1
;
CAXI4DMAOl01l
<=
{
{
(
CAXI4DMAl0OI
-
CAXI4DMAI1OI
)
{
1
'b
0
}
}
,
CAXI4DMAl1IIl
}
;
CAXI4DMAIO01l
<=
CAXI4DMAI1IIl
;
CAXI4DMAOI01l
<=
CAXI4DMAIIIIl
;
CAXI4DMAlI01l
<=
CAXI4DMAOIOIl
;
CAXI4DMAI1l0l
<=
CAXI4DMAlOOIl
;
CAXI4DMAOO1OI
<=
CAXI4DMAI000l
;
if
(
CAXI4DMAllllI
==
8
'b
00000001
)
begin
CAXI4DMAll01l
<=
PRI_0_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000010
)
begin
CAXI4DMAll01l
<=
PRI_1_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00000100
)
begin
CAXI4DMAll01l
<=
PRI_2_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00001000
)
begin
CAXI4DMAll01l
<=
PRI_3_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00010000
)
begin
CAXI4DMAll01l
<=
PRI_4_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
00100000
)
begin
CAXI4DMAll01l
<=
PRI_5_NUM_OF_BEATS
;
end
else
if
(
CAXI4DMAllllI
==
8
'b
01000000
)
begin
CAXI4DMAll01l
<=
PRI_6_NUM_OF_BEATS
;
end
else
begin
CAXI4DMAll01l
<=
PRI_7_NUM_OF_BEATS
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAOO10l
:
begin
if
(
CAXI4DMAOO1Ol
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAO101l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO10l
;
end
end
CAXI4DMAI101l
:
begin
if
(
CAXI4DMAlOlIl
)
begin
CAXI4DMAI0l1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAl101l
;
end
else
if
(
CAXI4DMAOIlIl
)
begin
CAXI4DMAO1l1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO11l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAI101l
;
end
end
CAXI4DMAI000l
:
begin
if
(
CAXI4DMAOOlIl
)
begin
CAXI4DMAlll1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO11l
;
end
else
if
(
CAXI4DMAIOlIl
)
begin
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO11l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAI000l
;
end
end
CAXI4DMAl101l
:
begin
if
(
CAXI4DMAlllIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAI0l1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAl101l
;
end
end
CAXI4DMAOO11l
:
begin
if
(
CAXI4DMAO0lIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAO1l1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO11l
;
end
end
CAXI4DMAIO11l
:
begin
if
(
CAXI4DMAOllIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAlll1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO11l
;
end
end
CAXI4DMAlO11l
:
begin
if
(
CAXI4DMAIllIl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO11l
;
end
end
CAXI4DMAOI11l
:
begin
if
(
CAXI4DMAIIlIl
)
begin
if
(
CAXI4DMAlIlIl
)
begin
CAXI4DMAl1l1l
<=
1
'b
1
;
CAXI4DMAO1Il
<=
1
'b
1
;
CAXI4DMAOl01l
<=
CAXI4DMAlIOIl
;
CAXI4DMAIO01l
<=
CAXI4DMAI1IIl
;
CAXI4DMAOI01l
<=
CAXI4DMAIIIIl
;
CAXI4DMAll01l
<=
PRI_0_NUM_OF_BEATS
;
CAXI4DMAOO1OI
<=
CAXI4DMAI101l
;
end
else
begin
CAXI4DMAI001l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAlOI
<=
1
'b
1
;
CAXI4DMAOII
<=
CAXI4DMAlI0OI
;
CAXI4DMAOO1OI
<=
CAXI4DMAOI11l
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIll1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAIll1l
<=
CAXI4DMAlll1l
;
end
end
assign
CAXI4DMAI0lIl
=
CAXI4DMAIll1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlO0ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAlO0ll
<=
CAXI4DMAOI0ll
;
end
end
assign
CAXI4DMAOllOI
=
CAXI4DMAlO0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO0l1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAO0l1l
<=
CAXI4DMAI0l1l
;
end
end
assign
CAXI4DMAl0lIl
=
CAXI4DMAO0l1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0l1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAl0l1l
<=
CAXI4DMAO1l1l
;
end
end
assign
CAXI4DMAO1lIl
=
CAXI4DMAl0l1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1l1l
<=
1
'b
0
;
end
else
begin
CAXI4DMAI1l1l
<=
CAXI4DMAl1l1l
;
end
end
assign
CAXI4DMAOI
=
CAXI4DMAI1l1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOO01l
<=
32
'b
0
;
end
else
begin
CAXI4DMAOO01l
<=
CAXI4DMAIO01l
;
end
end
assign
CAXI4DMAI101I
=
CAXI4DMAOO01l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlO01l
<=
2
'b
0
;
end
else
begin
CAXI4DMAlO01l
<=
CAXI4DMAOI01l
;
end
end
assign
CAXI4DMAl0
=
CAXI4DMAlO01l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAII01l
<=
3
'b
0
;
end
else
begin
CAXI4DMAII01l
<=
CAXI4DMAlI01l
;
end
end
assign
CAXI4DMAI1
=
CAXI4DMAII01l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO1l0l
<=
3
'b
0
;
end
else
begin
CAXI4DMAO1l0l
<=
CAXI4DMAI1l0l
;
end
end
assign
CAXI4DMAll
=
CAXI4DMAO1l0l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlI0Ol
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAlI0Ol
<=
CAXI4DMAOl01l
;
end
end
assign
CAXI4DMAlI0
=
CAXI4DMAlI0Ol
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIl01l
<=
{
CAXI4DMAI1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIl01l
<=
CAXI4DMAll01l
;
end
end
assign
CAXI4DMAIOI
=
CAXI4DMAIl01l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0Il
<=
1
'b
0
;
end
else
begin
CAXI4DMAl0Il
<=
CAXI4DMAO1Il
;
end
end
assign
CAXI4DMAI0
=
CAXI4DMAl0Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO001l
<=
1
'b
0
;
end
else
begin
CAXI4DMAO001l
<=
CAXI4DMAI001l
;
end
end
assign
CAXI4DMAl00Ol
=
CAXI4DMAO001l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl001l
<=
1
'b
0
;
end
else
begin
CAXI4DMAl001l
<=
CAXI4DMAO101l
;
end
end
assign
CAXI4DMAI10Ol
=
CAXI4DMAl001l
;
endmodule
