// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAOI11I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAO01lI
,
CAXI4DMAlI11I
,
CAXI4DMAOl11I
,
CAXI4DMAIlO0I
)
;
parameter
CAXI4DMAIl1lI
=
4
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAO01lI
;
input
CAXI4DMAlI11I
;
output
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAOl11I
;
output
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAIlO0I
;
localparam
[
1
:
0
]
CAXI4DMAO1OII
=
2
'b
01
;
localparam
[
1
:
0
]
CAXI4DMAOII1l
=
2
'b
10
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAO1O1l
;
reg
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAI1O1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAl1O1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAOOI1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAIOI1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAlOI1l
;
reg
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAIII1l
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAlII1l
;
reg
CAXI4DMAOlO0I
;
reg
CAXI4DMAOlI1l
;
reg
[
1
:
0
]
CAXI4DMAl10OI
;
reg
[
1
:
0
]
CAXI4DMAOO1OI
;
assign
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
1
:
0
]
&
CAXI4DMAI1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
assign
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
1
:
1
]
=
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
2
:
0
]
|
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
2
:
0
]
;
assign
CAXI4DMAl1O1l
[
0
]
=
1
'b
0
;
assign
CAXI4DMAOOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
&
~
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
assign
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
1
:
1
]
=
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
2
:
0
]
|
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
2
:
0
]
;
assign
CAXI4DMAIOI1l
[
0
]
=
1
'b
0
;
assign
CAXI4DMAlOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
1
:
0
]
&
~
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
assign
CAXI4DMAlII1l
[
CAXI4DMAIl1lI
-
1
:
0
]
=
(
|
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
)
?
CAXI4DMAOOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
:
CAXI4DMAlOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
CAXI4DMAIII1l
<=
{
CAXI4DMAIl1lI
{
1
'b
0
}
}
;
else
if
(
CAXI4DMAOlO0I
)
CAXI4DMAIII1l
<=
CAXI4DMAlII1l
;
else
if
(
CAXI4DMAOlI1l
)
CAXI4DMAIII1l
<=
{
CAXI4DMAIl1lI
{
1
'b
0
}
}
;
end
assign
CAXI4DMAIlO0I
=
CAXI4DMAIII1l
;
assign
CAXI4DMAOl11I
=
(
CAXI4DMAOlO0I
)
?
CAXI4DMAlII1l
:
{
CAXI4DMAIl1lI
{
1
'b
0
}
}
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1O1l
<=
{
CAXI4DMAIl1lI
{
1
'b
1
}
}
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
if
(
|
CAXI4DMAO1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
)
begin
CAXI4DMAI1O1l
<=
CAXI4DMAl1O1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
end
else
begin
CAXI4DMAI1O1l
<=
CAXI4DMAIOI1l
[
CAXI4DMAIl1lI
-
1
:
0
]
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAOlO0I
<=
1
'b
0
;
CAXI4DMAOlI1l
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
|
CAXI4DMAlII1l
)
begin
CAXI4DMAOlO0I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOII1l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAOII1l
:
begin
if
(
CAXI4DMAlI11I
)
begin
if
(
|
CAXI4DMAlII1l
)
begin
CAXI4DMAOlO0I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOII1l
;
end
else
begin
CAXI4DMAOlI1l
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOII1l
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
endmodule
