// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAllO1I
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAOlO1I
,
CAXI4DMAO1OOI
,
CAXI4DMAl11l
,
CAXI4DMAI0O1I
,
CAXI4DMAl0O1I
,
CAXI4DMAO1O1I
,
CAXI4DMAO1I0I
,
CAXI4DMAI1O1I
,
CAXI4DMAI011
,
CAXI4DMAI10
,
CAXI4DMAl1O1I
,
CAXI4DMAO10
,
CAXI4DMAl10
,
CAXI4DMAOOI1I
,
CAXI4DMAIOI1I
,
intDscrptrNum
,
CAXI4DMAlI0OI
,
CAXI4DMAO1IOI
,
CAXI4DMAlI1l
,
CAXI4DMAI1IlI
,
CAXI4DMAlOI1I
,
CAXI4DMAl1I0I
,
CAXI4DMAl010I
,
CAXI4DMAOII1I
,
CAXI4DMAIII1I
,
CAXI4DMAlII1I
,
CAXI4DMAOlI1I
,
CAXI4DMAIlI
,
CAXI4DMAllI
,
CAXI4DMAO0I
,
CAXI4DMAl0I
,
CAXI4DMAIlI1I
,
CAXI4DMAO1I
)
;
parameter
CAXI4DMAl1OI
=
133
;
parameter
CAXI4DMAl0OI
=
12
;
parameter
CAXI4DMAOIO1
=
2
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAOlO1I
;
input
CAXI4DMAO1OOI
;
input
[
31
:
0
]
CAXI4DMAl11l
;
input
CAXI4DMAI0O1I
;
input
CAXI4DMAl0O1I
;
input
CAXI4DMAO1O1I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO1I0I
;
input
[
31
:
0
]
CAXI4DMAI1O1I
;
input
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAI10
;
input
CAXI4DMAl10
;
input
CAXI4DMAl1O1I
;
input
[
1
:
0
]
CAXI4DMAO10
;
input
[
7
:
0
]
CAXI4DMAI011
;
output
reg
CAXI4DMAOOI1I
;
output
reg
CAXI4DMAIOI1I
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
intDscrptrNum
;
output
[
31
:
0
]
CAXI4DMAlI0OI
;
output
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAO1IOI
;
output
CAXI4DMAlI1l
;
output
CAXI4DMAI1IlI
;
output
CAXI4DMAlOI1I
;
output
CAXI4DMAl1I0I
;
output
reg
CAXI4DMAl010I
;
output
reg
CAXI4DMAOII1I
;
output
CAXI4DMAIII1I
;
output
reg
CAXI4DMAlII1I
;
output
reg
CAXI4DMAOlI1I
;
output
reg
CAXI4DMAIlI
;
output
reg
CAXI4DMAllI
;
output
reg
CAXI4DMAO0I
;
output
reg
CAXI4DMAl0I
;
output
reg
[
31
:
0
]
CAXI4DMAIlI1I
;
output
reg
[
7
:
0
]
CAXI4DMAO1I
;
localparam
[
7
:
0
]
CAXI4DMAO1OII
=
8
'b
00000001
;
localparam
[
7
:
0
]
CAXI4DMAl10Il
=
8
'b
00000010
;
localparam
[
7
:
0
]
CAXI4DMAOO1Il
=
8
'b
00000100
;
localparam
[
7
:
0
]
CAXI4DMAIO1Il
=
8
'b
00001000
;
localparam
[
7
:
0
]
CAXI4DMAlO1Il
=
8
'b
00010000
;
localparam
[
7
:
0
]
CAXI4DMAOI1Il
=
8
'b
00100000
;
localparam
[
7
:
0
]
CAXI4DMAII1Il
=
8
'b
01000000
;
localparam
[
7
:
0
]
CAXI4DMAlI1Il
=
8
'b
10000000
;
localparam
CAXI4DMAOl1Il
=
1
;
reg
[
7
:
0
]
CAXI4DMAl10OI
;
reg
[
7
:
0
]
CAXI4DMAOO1OI
;
reg
CAXI4DMAIl1Il
;
reg
CAXI4DMAll1Il
;
reg
CAXI4DMAO01Il
;
reg
CAXI4DMAI01Il
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl01Il
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO11Il
;
reg
[
31
:
0
]
CAXI4DMAI11Il
;
reg
[
31
:
0
]
CAXI4DMAl11Il
;
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAOOOll
;
reg
[
CAXI4DMAl1OI
-
1
:
0
]
CAXI4DMAIOOll
;
reg
CAXI4DMAO10II
;
reg
CAXI4DMAlOOll
;
reg
CAXI4DMAOIOll
;
reg
CAXI4DMAIIOll
;
reg
CAXI4DMAlIOll
;
reg
CAXI4DMAOlOll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAll1Il
<=
1
'b
0
;
CAXI4DMAI01Il
<=
CAXI4DMAO01Il
;
CAXI4DMAO11Il
<=
CAXI4DMAl01Il
;
CAXI4DMAl11Il
<=
CAXI4DMAI11Il
;
CAXI4DMAIOOll
<=
CAXI4DMAOOOll
;
CAXI4DMAlOOll
<=
CAXI4DMAO10II
;
CAXI4DMAIlI
<=
1
'b
0
;
CAXI4DMAllI
<=
1
'b
0
;
CAXI4DMAO0I
<=
1
'b
0
;
CAXI4DMAIlI1I
<=
32
'b
0
;
CAXI4DMAl0I
<=
1
'b
0
;
CAXI4DMAOlOll
<=
1
'b
0
;
CAXI4DMAOII1I
<=
1
'b
0
;
CAXI4DMAlII1I
<=
1
'b
0
;
CAXI4DMAOOI1I
<=
1
'b
0
;
CAXI4DMAIOI1I
<=
1
'b
0
;
CAXI4DMAIIOll
<=
1
'b
0
;
CAXI4DMAOlI1I
<=
1
'b
0
;
CAXI4DMAO1I
<=
8
'b
0
;
CAXI4DMAl010I
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAI0O1I
)
begin
CAXI4DMAllI
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10Il
;
end
else
if
(
CAXI4DMAO1O1I
)
begin
CAXI4DMAO0I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
+
CAXI4DMAOl1Il
;
CAXI4DMAOO1OI
<=
CAXI4DMAIO1Il
;
end
else
if
(
CAXI4DMAl0O1I
)
begin
CAXI4DMAO1I
<=
CAXI4DMAI011
;
CAXI4DMAl0I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
+
CAXI4DMAOl1Il
;
CAXI4DMAOO1OI
<=
CAXI4DMAOI1Il
;
end
else
if
(
CAXI4DMAO1OOI
)
begin
CAXI4DMAIlI
<=
1
'b
1
;
CAXI4DMAl010I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAl11l
;
CAXI4DMAOO1OI
<=
CAXI4DMAII1Il
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl10OI
;
end
end
CAXI4DMAl10Il
:
begin
if
(
CAXI4DMAl1O1I
)
begin
CAXI4DMAll1Il
<=
1
'b
1
;
CAXI4DMAI01Il
<=
&
CAXI4DMAO10
[
1
:
0
]
;
CAXI4DMAO11Il
<=
CAXI4DMAO1I0I
;
CAXI4DMAl11Il
<=
CAXI4DMAI1O1I
;
CAXI4DMAIOOll
<=
{
CAXI4DMAI10
[
133
:
14
]
,
&
CAXI4DMAO10
[
1
:
0
]
,
CAXI4DMAI10
[
12
:
0
]
}
;
CAXI4DMAlOOll
<=
CAXI4DMAl10
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO1Il
;
end
else
begin
CAXI4DMAllI
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10OI
;
end
end
CAXI4DMAOO1Il
:
begin
if
(
CAXI4DMAOlO1I
)
begin
CAXI4DMAI01Il
<=
1
'b
0
;
CAXI4DMAO11Il
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAl11Il
<=
32
'b
0
;
CAXI4DMAIOOll
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
CAXI4DMAlOOll
<=
1
'b
0
;
CAXI4DMAOII1I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAll1Il
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAOO1Il
;
end
end
CAXI4DMAIO1Il
:
begin
if
(
CAXI4DMAl1O1I
)
begin
CAXI4DMAlII1I
<=
1
'b
1
;
CAXI4DMAOlI1I
<=
&
CAXI4DMAO10
[
1
:
0
]
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAO0I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
+
CAXI4DMAOl1Il
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10OI
;
end
end
CAXI4DMAOI1Il
:
begin
if
(
CAXI4DMAl1O1I
)
begin
CAXI4DMAIIOll
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAlO1Il
;
end
else
begin
CAXI4DMAO1I
<=
CAXI4DMAI011
;
CAXI4DMAl0I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
+
CAXI4DMAOl1Il
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10OI
;
end
end
CAXI4DMAlO1Il
:
begin
if
(
CAXI4DMAI0O1I
)
begin
CAXI4DMAllI
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAI1O1I
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10Il
;
end
else
if
(
CAXI4DMAO1OOI
)
begin
CAXI4DMAIlI
<=
1
'b
1
;
CAXI4DMAl010I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAl11l
;
CAXI4DMAOO1OI
<=
CAXI4DMAII1Il
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAII1Il
:
begin
if
(
CAXI4DMAl1O1I
)
begin
CAXI4DMAll1Il
<=
1
'b
1
;
CAXI4DMAOlOll
<=
1
'b
1
;
CAXI4DMAI01Il
<=
CAXI4DMAO10
[
0
]
;
CAXI4DMAO11Il
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAl11Il
<=
CAXI4DMAl11l
;
CAXI4DMAIOOll
<=
CAXI4DMAI10
;
CAXI4DMAlOOll
<=
CAXI4DMAl10
;
CAXI4DMAOO1OI
<=
CAXI4DMAlI1Il
;
end
else
begin
CAXI4DMAIlI
<=
1
'b
1
;
CAXI4DMAl010I
<=
1
'b
1
;
CAXI4DMAIlI1I
<=
CAXI4DMAl11l
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10OI
;
end
end
CAXI4DMAlI1Il
:
begin
if
(
CAXI4DMAOlO1I
)
begin
CAXI4DMAI01Il
<=
1
'b
0
;
CAXI4DMAO11Il
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAl11Il
<=
32
'b
0
;
CAXI4DMAIOOll
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
CAXI4DMAlOOll
<=
1
'b
0
;
CAXI4DMAOOI1I
<=
1
'b
1
;
CAXI4DMAIOI1I
<=
CAXI4DMAO10II
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAll1Il
<=
1
'b
1
;
CAXI4DMAOlOll
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAl10OI
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIl1Il
<=
1
'b
0
;
end
else
begin
CAXI4DMAIl1Il
<=
CAXI4DMAll1Il
;
end
end
assign
CAXI4DMAl1I0I
=
CAXI4DMAIl1Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO01Il
<=
1
'b
0
;
end
else
begin
CAXI4DMAO01Il
<=
CAXI4DMAI01Il
;
end
end
assign
CAXI4DMAI1IlI
=
CAXI4DMAO01Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl01Il
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAl01Il
<=
CAXI4DMAO11Il
;
end
end
assign
intDscrptrNum
=
CAXI4DMAl01Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI11Il
<=
32
'b
0
;
end
else
begin
CAXI4DMAI11Il
<=
CAXI4DMAl11Il
;
end
end
assign
CAXI4DMAlI0OI
=
CAXI4DMAI11Il
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOOOll
<=
{
CAXI4DMAl1OI
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAOOOll
<=
CAXI4DMAIOOll
;
end
end
assign
CAXI4DMAO1IOI
=
CAXI4DMAOOOll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO10II
<=
1
'b
0
;
end
else
begin
CAXI4DMAO10II
<=
CAXI4DMAlOOll
;
end
end
assign
CAXI4DMAlI1l
=
CAXI4DMAO10II
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIOll
<=
1
'b
0
;
end
else
begin
CAXI4DMAOIOll
<=
CAXI4DMAIIOll
;
end
end
assign
CAXI4DMAIII1I
=
CAXI4DMAOIOll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlIOll
<=
1
'b
0
;
end
else
begin
CAXI4DMAlIOll
<=
CAXI4DMAOlOll
;
end
end
assign
CAXI4DMAlOI1I
=
CAXI4DMAlIOll
;
endmodule
