// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAI1OlI
(
CAXI4DMAI
,
CAXI4DMAOO1
,
CAXI4DMAIO1
,
CAXI4DMAlO1
,
CAXI4DMAIO1l
,
CAXI4DMAlI1
,
CAXI4DMAI1Il
)
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl1OlI
=
1
;
input
CAXI4DMAI
;
input
CAXI4DMAOO1
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIO1
;
input
[
31
:
0
]
CAXI4DMAlO1
;
input
CAXI4DMAIO1l
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlI1
;
output
[
31
:
0
]
CAXI4DMAI1Il
;
wire
[
19
:
0
]
CAXI4DMAl0I0l
;
wire
[
19
:
0
]
CAXI4DMAO1I0l
;
wire
CAXI4DMAI1I0l
;
assign
CAXI4DMAI1Il
=
{
CAXI4DMAl0I0l
[
11
:
0
]
,
CAXI4DMAO1I0l
[
19
:
0
]
}
;
assign
CAXI4DMAI1I0l
=
(
CAXI4DMAl1OlI
==
1
)
?
1
'b
0
:
1
'b
1
;
RAM1K20
CAXI4DMAl1I0l
(
.A_DOUT
(
CAXI4DMAl0I0l
)
,
.B_DOUT
(
CAXI4DMAO1I0l
)
,
.DB_DETECT
(
)
,
.SB_CORRECT
(
)
,
.ACCESS_BUSY
(
)
,
.A_ADDR
(
{
{
(
9
-
CAXI4DMAOIO1
)
{
1
'b
1
}
}
,
CAXI4DMAlI1
[
CAXI4DMAOIO1
-
1
:
0
]
,
{
5
{
1
'b
0
}
}
}
)
,
.A_BLK_EN
(
3
'b
111
)
,
.A_CLK
(
CAXI4DMAI
)
,
.A_DIN
(
{
{
8
{
1
'b
0
}
}
,
CAXI4DMAlO1
[
31
:
20
]
}
)
,
.A_REN
(
CAXI4DMAIO1l
)
,
.A_WEN
(
2
'b
11
)
,
.A_DOUT_EN
(
1
'b
1
)
,
.A_DOUT_ARST_N
(
1
'b
1
)
,
.A_DOUT_SRST_N
(
1
'b
1
)
,
.B_ADDR
(
{
{
(
9
-
CAXI4DMAOIO1
)
{
1
'b
1
}
}
,
CAXI4DMAIO1
[
CAXI4DMAOIO1
-
1
:
0
]
,
{
5
{
1
'b
0
}
}
}
)
,
.B_BLK_EN
(
{
CAXI4DMAOO1
,
2
'b
11
}
)
,
.B_CLK
(
CAXI4DMAI
)
,
.B_DIN
(
{
CAXI4DMAlO1
[
19
:
0
]
}
)
,
.B_REN
(
1
'b
1
)
,
.B_WEN
(
2
'b
11
)
,
.B_DOUT_EN
(
1
'b
1
)
,
.B_DOUT_ARST_N
(
1
'b
1
)
,
.B_DOUT_SRST_N
(
1
'b
1
)
,
.ECC_EN
(
1
'b
0
)
,
.BUSY_FB
(
1
'b
0
)
,
.A_WIDTH
(
3
'b
101
)
,
.A_WMODE
(
2
'b
00
)
,
.A_BYPASS
(
CAXI4DMAI1I0l
)
,
.B_WIDTH
(
3
'b
101
)
,
.B_WMODE
(
2
'b
00
)
,
.B_BYPASS
(
CAXI4DMAI1I0l
)
,
.ECC_BYPASS
(
1
'b
0
)
)
;
endmodule
