// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28871 $
// SVN $Date: 2017-02-13 03:32:54 +0000 (Mon, 13 Feb 2017) $
module
CAXI4DMAlO1Ol
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAO011I
,
CAXI4DMAI011I
,
CAXI4DMAl011I
,
CAXI4DMAO111I
,
CAXI4DMAI111I
,
CAXI4DMAII1Ol
,
CAXI4DMAIOOOl
,
CAXI4DMAI1lOl
,
CAXI4DMAOI0Ol
,
CAXI4DMAO1lOl
,
CAXI4DMAl0lOl
,
CAXI4DMAIIlOl
,
CAXI4DMAlOOOl
,
CAXI4DMAI0IOl
,
CAXI4DMAl111I
,
CAXI4DMAOOOOl
,
CAXI4DMAOIOOl
,
CAXI4DMAIIOOl
,
CAXI4DMAlIOOl
,
CAXI4DMAIOlOl
,
CAXI4DMAlI0
,
CAXI4DMAOlOOl
,
CAXI4DMAIlOOl
,
CAXI4DMAllOOl
,
CAXI4DMAO0OOl
,
CAXI4DMAlI1Ol
,
CAXI4DMAI00
,
CAXI4DMAl00Ol
,
CAXI4DMAI0OOl
,
CAXI4DMAl0OOl
,
CAXI4DMAO1OOl
,
CAXI4DMAI10Ol
,
CAXI4DMAO10Ol
,
CAXI4DMAI1I1I
,
CAXI4DMAOII1I
,
CAXI4DMAIII1I
,
CAXI4DMAIO0lI
,
CAXI4DMAOlllI
,
CAXI4DMAI1OOl
,
CAXI4DMAl1OOl
,
CAXI4DMAOO10I
,
CAXI4DMAlIlOI
,
CAXI4DMAOllOI
,
CAXI4DMAIllOI
,
CAXI4DMAI1l0I
,
CAXI4DMAO010I
,
CAXI4DMAl1l0I
,
CAXI4DMAI010I
,
CAXI4DMAOOIOl
,
CAXI4DMAIOIOl
,
CAXI4DMAlOIOl
,
CAXI4DMAOIIOl
,
CAXI4DMAIII
,
CAXI4DMAlII
,
CAXI4DMAOlI
,
CAXI4DMAIIIOl
,
CAXI4DMAlIIOl
,
CAXI4DMAOlIOl
,
CAXI4DMAOO1Ol
,
CAXI4DMAl10Ol
,
CAXI4DMAI1l1
,
CAXI4DMAl1l1
,
CAXI4DMAOl1Ol
,
CAXI4DMAl0I
,
CAXI4DMAIl1Ol
,
CAXI4DMAll1Ol
,
CAXI4DMAO1I
,
CAXI4DMAl1lOl
,
CAXI4DMAOl1l
,
CAXI4DMAIl1l
)
;
parameter
NUM_INT_BDS
=
4
;
parameter
CAXI4DMAOIO1
=
2
;
parameter
CAXI4DMAl0OI
=
23
;
parameter
CAXI4DMAO1OI
=
12
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAO011I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI011I
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAl011I
;
input
[
31
:
0
]
CAXI4DMAO111I
;
input
CAXI4DMAI111I
;
input
CAXI4DMAl111I
;
input
CAXI4DMAO1lOl
;
input
[
31
:
0
]
CAXI4DMAII1Ol
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIOOOl
;
input
[
7
:
0
]
CAXI4DMAI1lOl
;
input
CAXI4DMAOI0Ol
;
input
CAXI4DMAl0lOl
;
input
[
1
:
0
]
CAXI4DMAIIlOl
;
input
CAXI4DMAlOOOl
;
input
CAXI4DMAI0IOl
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOIOOl
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIIOOl
;
input
[
31
:
0
]
CAXI4DMAlIOOl
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAIOlOl
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI0
;
input
CAXI4DMAOOOOl
;
input
CAXI4DMAOlOOl
;
input
CAXI4DMAIlOOl
;
input
CAXI4DMAllOOl
;
input
CAXI4DMAO0OOl
;
input
[
CAXI4DMAO1OI
-
1
:
0
]
CAXI4DMAlI1Ol
;
input
CAXI4DMAI00
;
input
CAXI4DMAl00Ol
;
input
CAXI4DMAI0OOl
;
input
CAXI4DMAl0OOl
;
input
CAXI4DMAO1OOl
;
input
CAXI4DMAI10Ol
;
input
CAXI4DMAO10Ol
;
input
CAXI4DMAI1I1I
;
input
CAXI4DMAOII1I
;
input
CAXI4DMAIII1I
;
output
reg
CAXI4DMAIO0lI
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOlllI
;
output
reg
[
1
:
0
]
CAXI4DMAI1OOl
;
output
reg
[
1
:
0
]
CAXI4DMAl1OOl
;
output
CAXI4DMAOO10I
;
output
CAXI4DMAlIlOI
;
output
CAXI4DMAOllOI
;
output
CAXI4DMAIllOI
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI1l0I
;
output
CAXI4DMAO010I
;
output
[
31
:
0
]
CAXI4DMAl1l0I
;
output
CAXI4DMAI010I
;
output
reg
CAXI4DMAOOIOl
;
output
reg
CAXI4DMAIOIOl
;
output
reg
CAXI4DMAlOIOl
;
output
reg
CAXI4DMAOIIOl
;
output
reg
CAXI4DMAIII
;
output
reg
[
31
:
0
]
CAXI4DMAlII
;
output
reg
[
1
:
0
]
CAXI4DMAOlI
;
output
reg
CAXI4DMAIIIOl
;
output
reg
CAXI4DMAlIIOl
;
output
reg
CAXI4DMAOlIOl
;
output
reg
CAXI4DMAOO1Ol
;
output
reg
CAXI4DMAl10Ol
;
output
reg
CAXI4DMAI1l1
;
output
reg
CAXI4DMAl1l1
;
output
CAXI4DMAOl1Ol
;
output
CAXI4DMAl0I
;
output
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIl1Ol
;
output
[
31
:
0
]
CAXI4DMAll1Ol
;
output
[
7
:
0
]
CAXI4DMAO1I
;
output
reg
CAXI4DMAl1lOl
;
output
CAXI4DMAOl1l
;
output
CAXI4DMAIl1l
;
reg
[
13
:
0
]
CAXI4DMAl10OI
;
reg
[
13
:
0
]
CAXI4DMAOO1OI
;
reg
CAXI4DMAl1Ill
;
reg
CAXI4DMAOOlll
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIOlll
[
0
:
1
]
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlOlll
[
0
:
1
]
;
reg
CAXI4DMAOIlll
;
reg
CAXI4DMAIIlll
;
reg
CAXI4DMAlIlll
;
reg
CAXI4DMAOllll
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIllll
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAlllll
;
reg
[
31
:
0
]
CAXI4DMAO0lll
;
reg
[
31
:
0
]
CAXI4DMAI0lll
;
reg
[
7
:
0
]
CAXI4DMAl0lll
;
reg
[
7
:
0
]
CAXI4DMAO1lll
;
reg
CAXI4DMAI1lll
;
reg
CAXI4DMAl1lll
;
reg
CAXI4DMAOO0ll
;
reg
CAXI4DMAIO0ll
;
reg
CAXI4DMAlO0ll
;
reg
CAXI4DMAOI0ll
;
reg
CAXI4DMAII0ll
;
reg
CAXI4DMAlI0ll
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAOl0ll
;
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAIl0ll
;
reg
CAXI4DMAll0ll
;
reg
CAXI4DMAO00ll
;
reg
[
31
:
0
]
CAXI4DMAI00ll
;
reg
[
31
:
0
]
CAXI4DMAl00ll
;
reg
CAXI4DMAO10ll
;
reg
CAXI4DMAI10ll
;
reg
CAXI4DMAl10ll
;
reg
CAXI4DMAOO1ll
;
reg
CAXI4DMAIO1ll
;
reg
CAXI4DMAlO1ll
;
reg
CAXI4DMAOI1ll
;
reg
[
31
:
0
]
CAXI4DMAII1ll
;
reg
[
1
:
0
]
CAXI4DMAlI1ll
;
localparam
[
13
:
0
]
CAXI4DMAO1OII
=
14
'b
00000000000001
;
localparam
[
13
:
0
]
CAXI4DMAOl1ll
=
14
'b
00000000000010
;
localparam
[
13
:
0
]
CAXI4DMAIl1ll
=
14
'b
00000000000100
;
localparam
[
13
:
0
]
CAXI4DMAll1ll
=
14
'b
00000000001000
;
localparam
[
13
:
0
]
CAXI4DMAO01ll
=
14
'b
00000000010000
;
localparam
[
13
:
0
]
CAXI4DMAI01ll
=
14
'b
00000000100000
;
localparam
[
13
:
0
]
CAXI4DMAl01ll
=
14
'b
00000001000000
;
localparam
[
13
:
0
]
CAXI4DMAO11ll
=
14
'b
00000010000000
;
localparam
[
13
:
0
]
CAXI4DMAI11ll
=
14
'b
00000100000000
;
localparam
[
13
:
0
]
CAXI4DMAl11ll
=
14
'b
00001000000000
;
localparam
[
13
:
0
]
CAXI4DMAOOO0l
=
14
'b
00010000000000
;
localparam
[
13
:
0
]
CAXI4DMAIOO0l
=
14
'b
00100000000000
;
localparam
[
13
:
0
]
CAXI4DMAlOO0l
=
14
'b
01000000000000
;
localparam
[
13
:
0
]
CAXI4DMAOIO0l
=
14
'b
10000000000000
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1l1
<=
1
'b
0
;
end
else
begin
CAXI4DMAI1l1
<=
CAXI4DMAl1Ill
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl1l1
<=
1
'b
0
;
end
else
begin
CAXI4DMAl1l1
<=
CAXI4DMAOOlll
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIlll
<=
1
'b
0
;
end
else
begin
CAXI4DMAOIlll
<=
CAXI4DMAIIlll
;
end
end
assign
CAXI4DMAOl1Ol
=
CAXI4DMAOIlll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlIlll
<=
1
'b
0
;
end
else
begin
CAXI4DMAlIlll
<=
CAXI4DMAOllll
;
end
end
assign
CAXI4DMAl0I
=
CAXI4DMAlIlll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIllll
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAIllll
<=
CAXI4DMAlllll
;
end
end
assign
CAXI4DMAIl1Ol
=
CAXI4DMAIllll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO0lll
<=
32
'b
0
;
end
else
begin
CAXI4DMAO0lll
<=
CAXI4DMAI0lll
;
end
end
assign
CAXI4DMAll1Ol
=
CAXI4DMAO0lll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0lll
<=
8
'b
0
;
end
else
begin
CAXI4DMAl0lll
<=
CAXI4DMAO1lll
;
end
end
assign
CAXI4DMAO1I
=
CAXI4DMAl0lll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI1lll
<=
1
'b
0
;
end
else
begin
CAXI4DMAI1lll
<=
CAXI4DMAl1lll
;
end
end
assign
CAXI4DMAOO10I
=
CAXI4DMAI1lll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOO0ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAOO0ll
<=
CAXI4DMAIO0ll
;
end
end
assign
CAXI4DMAlIlOI
=
CAXI4DMAOO0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlO0ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAlO0ll
<=
CAXI4DMAOI0ll
;
end
end
assign
CAXI4DMAOllOI
=
CAXI4DMAlO0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAII0ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAII0ll
<=
CAXI4DMAlI0ll
;
end
end
assign
CAXI4DMAIllOI
=
CAXI4DMAII0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOl0ll
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
end
else
begin
CAXI4DMAOl0ll
<=
CAXI4DMAIl0ll
;
end
end
assign
CAXI4DMAI1l0I
=
CAXI4DMAOl0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAll0ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAll0ll
<=
CAXI4DMAO00ll
;
end
end
assign
CAXI4DMAO010I
=
CAXI4DMAll0ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI00ll
<=
32
'b
0
;
end
else
begin
CAXI4DMAI00ll
<=
CAXI4DMAl00ll
;
end
end
assign
CAXI4DMAl1l0I
=
CAXI4DMAI00ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO10ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAO10ll
<=
CAXI4DMAI10ll
;
end
end
assign
CAXI4DMAI010I
=
CAXI4DMAO10ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAl10ll
<=
CAXI4DMAOO1ll
;
end
end
assign
CAXI4DMAOl1l
=
CAXI4DMAl10ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO1ll
<=
1
'b
0
;
end
else
begin
CAXI4DMAIO1ll
<=
CAXI4DMAlO1ll
;
end
end
assign
CAXI4DMAIl1l
=
CAXI4DMAIO1ll
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIII
<=
1
'b
0
;
end
else
begin
CAXI4DMAIII
<=
CAXI4DMAOI1ll
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAlII
<=
32
'b
0
;
end
else
begin
CAXI4DMAlII
<=
CAXI4DMAII1ll
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOlI
<=
2
'b
0
;
end
else
begin
CAXI4DMAOlI
<=
CAXI4DMAlI1ll
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAIOlll
[
0
]
=
CAXI4DMAI011I
;
CAXI4DMAIOlll
[
1
]
=
CAXI4DMAl011I
;
CAXI4DMAlOlll
[
0
]
=
CAXI4DMAOIOOl
;
CAXI4DMAlOlll
[
1
]
=
CAXI4DMAIIOOl
;
end
always
@
(
*
)
begin
CAXI4DMAI1OOl
[
0
]
<=
1
'b
0
;
CAXI4DMAI1OOl
[
1
]
<=
1
'b
0
;
CAXI4DMAOOIOl
<=
1
'b
0
;
CAXI4DMAIOIOl
<=
1
'b
0
;
CAXI4DMAlOIOl
<=
1
'b
0
;
CAXI4DMAOIIOl
<=
1
'b
0
;
CAXI4DMAl1Ill
<=
CAXI4DMAI1l1
;
CAXI4DMAl1lll
<=
1
'b
0
;
CAXI4DMAIO0ll
<=
1
'b
0
;
CAXI4DMAOI0ll
<=
1
'b
0
;
CAXI4DMAlI0ll
<=
1
'b
0
;
CAXI4DMAIl0ll
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAO00ll
<=
1
'b
0
;
CAXI4DMAl00ll
<=
32
'b
0
;
CAXI4DMAl1OOl
[
0
]
<=
1
'b
0
;
CAXI4DMAl1OOl
[
1
]
<=
1
'b
0
;
CAXI4DMAIIIOl
<=
1
'b
0
;
CAXI4DMAlIIOl
<=
1
'b
0
;
CAXI4DMAOOlll
<=
CAXI4DMAl1l1
;
CAXI4DMAIO0lI
<=
1
'b
0
;
CAXI4DMAOlllI
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAIIlll
<=
1
'b
0
;
CAXI4DMAlllll
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAI0lll
<=
32
'b
0
;
CAXI4DMAOlIOl
<=
1
'b
0
;
CAXI4DMAOllll
<=
1
'b
0
;
CAXI4DMAO1lll
<=
8
'b
0
;
CAXI4DMAl1lOl
<=
1
'b
0
;
CAXI4DMAI10ll
<=
1
'b
0
;
CAXI4DMAOO1ll
<=
1
'b
0
;
CAXI4DMAlO1ll
<=
1
'b
0
;
CAXI4DMAOI1ll
<=
1
'b
0
;
CAXI4DMAII1ll
<=
32
'b
0
;
CAXI4DMAlI1ll
<=
2
'b
0
;
CAXI4DMAOO1Ol
<=
1
'b
0
;
CAXI4DMAl10Ol
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAO1OII
:
begin
if
(
CAXI4DMAI10Ol
)
begin
if
(
CAXI4DMAl0lOl
)
begin
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAIIlll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAII1Ol
;
CAXI4DMAOO1OI
<=
CAXI4DMAl11ll
;
end
else
begin
CAXI4DMAl1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOO1Ol
<=
1
'b
1
;
CAXI4DMAl10Ol
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAl1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOO1Ol
<=
1
'b
1
;
CAXI4DMAl10Ol
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
if
(
CAXI4DMAO1OOl
)
begin
CAXI4DMAI1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAOlIOl
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
if
(
CAXI4DMAl00Ol
)
begin
CAXI4DMAI1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
if
(
CAXI4DMAl0OOl
)
begin
CAXI4DMAIO0lI
<=
1
'b
1
;
CAXI4DMAOlllI
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
if
(
CAXI4DMAI1l1
==
CAXI4DMAl1l1
)
begin
if
(
!
CAXI4DMAO011I
)
begin
if
(
CAXI4DMAIOlll
[
!
CAXI4DMAI1l1
]
==
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
)
begin
CAXI4DMAI1OOl
[
!
CAXI4DMAI1l1
]
<=
1
'b
1
;
end
end
CAXI4DMAOO1OI
<=
CAXI4DMAOl1ll
;
end
else
begin
if
(
!
CAXI4DMAO011I
)
begin
if
(
CAXI4DMAIOlll
[
!
CAXI4DMAI1l1
]
==
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
)
begin
CAXI4DMAI1OOl
[
!
CAXI4DMAI1l1
]
<=
1
'b
1
;
end
end
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI0IOl
;
CAXI4DMAl00ll
<=
CAXI4DMAlIOOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAIl1ll
;
end
end
else
if
(
CAXI4DMAIlOOl
)
begin
CAXI4DMAIO0lI
<=
1
'b
1
;
CAXI4DMAOlllI
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
if
(
!
CAXI4DMAlOOOl
)
begin
if
(
CAXI4DMAlOlll
[
!
CAXI4DMAl1l1
]
==
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
)
begin
CAXI4DMAl1OOl
[
!
CAXI4DMAl1l1
]
<=
1
'b
1
;
end
end
if
(
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
==
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAI01ll
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAl01ll
;
end
end
else
if
(
CAXI4DMAOlOOl
)
begin
if
(
CAXI4DMAIOOOl
==
{
{
(
CAXI4DMAl0OI
-
CAXI4DMAO1OI
)
{
1
'b
0
}
}
,
CAXI4DMAlI1Ol
}
)
begin
if
(
CAXI4DMAI111I
)
begin
CAXI4DMAOllll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAO111I
;
CAXI4DMAO1lll
<=
CAXI4DMAI1lOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAI11ll
;
end
else
begin
if
(
CAXI4DMAl0lOl
)
begin
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAIIlll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAII1Ol
;
end
if
(
CAXI4DMAOI0Ol
)
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOOO0l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO11ll
;
end
end
else
begin
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl11ll
;
end
else
begin
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAO11ll
;
end
end
end
else
begin
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
if
(
CAXI4DMAI0OOl
)
begin
if
(
CAXI4DMAIOlOl
==
{
{
(
CAXI4DMAl0OI
-
CAXI4DMAO1OI
)
{
1
'b
0
}
}
,
CAXI4DMAlI0
}
)
begin
if
(
CAXI4DMAl111I
)
begin
if
(
CAXI4DMAOOOOl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
if
(
CAXI4DMAO0OOl
||
CAXI4DMAllOOl
)
begin
CAXI4DMAOI1ll
<=
1
'b
1
;
CAXI4DMAII1ll
<=
CAXI4DMAO111I
;
CAXI4DMAlI1ll
<=
CAXI4DMAIIlOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAOIO0l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
CAXI4DMAI11ll
:
begin
if
(
CAXI4DMAIII1I
)
begin
if
(
CAXI4DMAl0lOl
)
begin
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAIIlll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAII1Ol
;
end
if
(
CAXI4DMAOI0Ol
)
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOOO0l
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO11ll
;
end
end
else
begin
if
(
CAXI4DMAO1lOl
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAl11ll
;
end
else
begin
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAO11ll
;
end
end
else
begin
CAXI4DMAOllll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAO111I
;
CAXI4DMAO1lll
<=
CAXI4DMAI1lOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAI11ll
;
end
end
CAXI4DMAO11ll
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAO11ll
;
end
end
CAXI4DMAl11ll
:
begin
if
(
CAXI4DMAOII1I
)
begin
if
(
CAXI4DMAI10Ol
)
begin
CAXI4DMAl1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOO1Ol
<=
1
'b
1
;
CAXI4DMAl10Ol
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
end
else
begin
CAXI4DMAIIlll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAII1Ol
;
CAXI4DMAOO1OI
<=
CAXI4DMAl11ll
;
end
end
CAXI4DMAOOO0l
:
begin
if
(
CAXI4DMAI1I1I
)
begin
if
(
CAXI4DMAOII1I
)
begin
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAIIlll
<=
1
'b
1
;
CAXI4DMAlllll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI0lll
<=
CAXI4DMAII1Ol
;
CAXI4DMAOO1OI
<=
CAXI4DMAl11ll
;
end
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
if
(
CAXI4DMAOII1I
)
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO11ll
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOOO0l
;
end
end
end
CAXI4DMAI01ll
:
begin
if
(
CAXI4DMAl0OOl
|
CAXI4DMAI0OOl
)
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
if
(
CAXI4DMAl0OOl
)
begin
CAXI4DMAlIIOl
<=
1
'b
1
;
end
else
begin
CAXI4DMAIIIOl
<=
1
'b
1
;
end
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAl01ll
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAI01ll
;
end
end
CAXI4DMAl01ll
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAIOIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI111I
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAl01ll
;
end
end
CAXI4DMAIl1ll
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAlIIOl
<=
1
'b
1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI0IOl
;
CAXI4DMAl00ll
<=
CAXI4DMAlIOOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAIl1ll
;
end
end
CAXI4DMAOl1ll
:
begin
if
(
CAXI4DMAIlOOl
)
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI0IOl
;
CAXI4DMAl00ll
<=
CAXI4DMAlIOOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAll1ll
;
end
else
if
(
CAXI4DMAOlOOl
)
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI0IOl
;
CAXI4DMAl00ll
<=
CAXI4DMAlIOOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAO01ll
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAOl1ll
;
end
end
CAXI4DMAll1ll
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAIOIOl
<=
1
'b
1
;
CAXI4DMAlIIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI0IOl
;
CAXI4DMAl00ll
<=
CAXI4DMAlIOOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAll1ll
;
end
end
CAXI4DMAO01ll
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAl1lOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAl1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAOOIOl
<=
1
'b
1
;
CAXI4DMAlIIOl
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAlI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAlOlll
[
CAXI4DMAl1l1
]
;
CAXI4DMAO00ll
<=
CAXI4DMAI0IOl
;
CAXI4DMAl00ll
<=
CAXI4DMAlIOOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAO01ll
;
end
end
CAXI4DMAlOO0l
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAlOIOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAl1l1
]
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI10ll
<=
1
'b
1
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAlOO0l
;
end
end
CAXI4DMAIOO0l
:
begin
if
(
CAXI4DMAI1I1I
)
begin
CAXI4DMAOIIOl
<=
1
'b
1
;
CAXI4DMAI1OOl
[
CAXI4DMAI1l1
]
<=
1
'b
1
;
CAXI4DMAl1Ill
<=
~
CAXI4DMAI1l1
;
CAXI4DMAOOlll
<=
~
CAXI4DMAl1l1
;
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
else
begin
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI10ll
<=
1
'b
1
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAIOO0l
;
end
end
CAXI4DMAOIO0l
:
begin
if
(
CAXI4DMAI00
)
begin
if
(
CAXI4DMAO0OOl
)
begin
CAXI4DMAlO1ll
<=
1
'b
1
;
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAOI0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI10ll
<=
1
'b
1
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAIOO0l
;
end
else
begin
CAXI4DMAOO1ll
<=
1
'b
1
;
CAXI4DMAl1lll
<=
1
'b
1
;
CAXI4DMAIO0ll
<=
1
'b
1
;
CAXI4DMAIl0ll
<=
CAXI4DMAIOlll
[
CAXI4DMAI1l1
]
;
CAXI4DMAI10ll
<=
1
'b
1
;
CAXI4DMAl00ll
<=
CAXI4DMAO111I
;
CAXI4DMAOO1OI
<=
CAXI4DMAlOO0l
;
end
end
else
begin
CAXI4DMAOI1ll
<=
1
'b
1
;
CAXI4DMAII1ll
<=
CAXI4DMAO111I
;
CAXI4DMAlI1ll
<=
CAXI4DMAIIlOl
;
CAXI4DMAOO1OI
<=
CAXI4DMAOIO0l
;
end
end
default
:
begin
CAXI4DMAOO1OI
<=
CAXI4DMAO1OII
;
end
endcase
end
endmodule
