// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAII1lI
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAO01lI
,
CAXI4DMAlO0lI
,
CAXI4DMAIO0lI
,
CAXI4DMAO00lI
,
CAXI4DMAI01lI
,
CAXI4DMAl01lI
,
CAXI4DMAO11lI
,
CAXI4DMAI11lI
,
CAXI4DMAl11lI
,
CAXI4DMAOOO0I
,
CAXI4DMAIOO0I
,
CAXI4DMAlOO0I
,
CAXI4DMAOO0lI
,
CAXI4DMAOIO0I
,
strDscrptr
,
intDscrptrNum
,
CAXI4DMAllllI
)
;
parameter
CAXI4DMAlI1lI
=
4
;
parameter
CAXI4DMAOl1lI
=
2
;
parameter
CAXI4DMAIl1lI
=
4
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAO01lI
;
input
CAXI4DMAlO0lI
;
input
CAXI4DMAIO0lI
;
input
CAXI4DMAO00lI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAI01lI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAl01lI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAO11lI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAI11lI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAl11lI
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAOOO0I
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAIOO0I
;
input
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAlOO0I
;
output
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAOO0lI
;
output
reg
CAXI4DMAOIO0I
;
output
reg
strDscrptr
;
output
reg
[
CAXI4DMAOl1lI
-
1
:
0
]
intDscrptrNum
;
output
reg
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAllllI
;
localparam
CAXI4DMAIlOll
=
0
;
localparam
CAXI4DMAllOll
=
1
;
reg
CAXI4DMAl10OI
;
reg
CAXI4DMAOO1OI
;
reg
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAO0Oll
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAI0Oll
;
reg
CAXI4DMAOlO0I
;
wire
[
CAXI4DMAOl1lI
-
1
:
0
]
CAXI4DMAl0Oll
;
wire
CAXI4DMAO1Oll
;
wire
[
CAXI4DMAIl1lI
-
1
:
0
]
CAXI4DMAI1Oll
;
generate
if
(
CAXI4DMAIl1lI
==
1
)
begin
assign
CAXI4DMAI0Oll
=
CAXI4DMAO01lI
;
end
else
if
(
CAXI4DMAIl1lI
>
1
)
begin
assign
CAXI4DMAI1Oll
[
CAXI4DMAIl1lI
-
1
:
1
]
=
CAXI4DMAI1Oll
[
CAXI4DMAIl1lI
-
2
:
0
]
|
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
2
:
0
]
;
assign
CAXI4DMAI1Oll
[
0
]
=
1
'b
0
;
assign
CAXI4DMAI0Oll
[
CAXI4DMAIl1lI
-
1
:
0
]
=
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
1
:
0
]
&
~
CAXI4DMAI1Oll
[
CAXI4DMAIl1lI
-
1
:
0
]
;
end
endgenerate
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO0Oll
<=
{
CAXI4DMAIl1lI
{
1
'b
0
}
}
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
CAXI4DMAO0Oll
<=
CAXI4DMAI0Oll
;
end
end
assign
CAXI4DMAOO0lI
[
CAXI4DMAIl1lI
-
1
:
0
]
=
(
CAXI4DMAOlO0I
)
?
CAXI4DMAI0Oll
[
CAXI4DMAIl1lI
-
1
:
0
]
:
{
CAXI4DMAIl1lI
{
1
'b
0
}
}
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAOIO0I
<=
1
'b
0
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
CAXI4DMAOIO0I
<=
1
'b
1
;
end
else
if
(
CAXI4DMAIO0lI
)
begin
CAXI4DMAOIO0I
<=
1
'b
0
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAllllI
<=
{
CAXI4DMAIl1lI
{
1
'b
0
}
}
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
CAXI4DMAllllI
<=
CAXI4DMAI0Oll
[
CAXI4DMAIl1lI
-
1
:
0
]
;
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
intDscrptrNum
<=
{
CAXI4DMAOl1lI
{
1
'b
0
}
}
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
intDscrptrNum
<=
CAXI4DMAl0Oll
;
end
end
assign
CAXI4DMAl0Oll
=
(
CAXI4DMAI0Oll
==
8
'b
00000010
)
?
CAXI4DMAl01lI
:
(
CAXI4DMAI0Oll
==
8
'b
00000100
)
?
CAXI4DMAO11lI
:
(
CAXI4DMAI0Oll
==
8
'b
00001000
)
?
CAXI4DMAI11lI
:
(
CAXI4DMAI0Oll
==
8
'b
00010000
)
?
CAXI4DMAl11lI
:
(
CAXI4DMAI0Oll
==
8
'b
00100000
)
?
CAXI4DMAOOO0I
:
(
CAXI4DMAI0Oll
==
8
'b
01000000
)
?
CAXI4DMAIOO0I
:
(
CAXI4DMAI0Oll
==
8
'b
10000000
)
?
CAXI4DMAlOO0I
:
CAXI4DMAI01lI
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
strDscrptr
<=
1
'b
0
;
end
else
if
(
CAXI4DMAOlO0I
)
begin
strDscrptr
<=
CAXI4DMAO1Oll
;
end
end
assign
CAXI4DMAO1Oll
=
(
CAXI4DMAI0Oll
==
8
'b
00000001
)
?
CAXI4DMAO00lI
:
1
'b
0
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl10OI
<=
CAXI4DMAIlOll
;
end
else
begin
CAXI4DMAl10OI
<=
CAXI4DMAOO1OI
;
end
end
always
@
(
*
)
begin
CAXI4DMAOlO0I
<=
1
'b
0
;
case
(
CAXI4DMAl10OI
)
CAXI4DMAIlOll
:
begin
if
(
|
CAXI4DMAO01lI
[
CAXI4DMAIl1lI
-
1
:
0
]
)
begin
CAXI4DMAOlO0I
<=
1
'b
1
;
CAXI4DMAOO1OI
<=
CAXI4DMAllOll
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIlOll
;
end
end
CAXI4DMAllOll
:
begin
if
(
CAXI4DMAlO0lI
)
begin
CAXI4DMAOO1OI
<=
CAXI4DMAIlOll
;
end
else
begin
CAXI4DMAOO1OI
<=
CAXI4DMAllOll
;
end
end
endcase
end
endmodule
