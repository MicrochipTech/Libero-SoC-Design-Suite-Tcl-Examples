// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// SVN Revision Information:
// SVN $Revision: 28772 $
// SVN $Date: 2017-02-09 20:06:50 +0000 (Thu, 09 Feb 2017) $
module
CAXI4DMAO01Ol
(
CAXI4DMAI
,
CAXI4DMAl
,
CAXI4DMAIlllI
,
CAXI4DMAI0llI
,
CAXI4DMAOIl1I
,
CAXI4DMAlOl1I
,
CAXI4DMAIIl1I
,
CAXI4DMAOll1I
,
CAXI4DMAIll1I
,
CAXI4DMAlll1I
,
CAXI4DMAOO01I
,
CAXI4DMAO0l1I
,
CAXI4DMAl100I
,
CAXI4DMAI0l1I
,
CAXI4DMAl0l1I
,
CAXI4DMAO1l1I
,
CAXI4DMAl01Ol
,
CAXI4DMAl1OOl
,
CAXI4DMAl1l1
,
CAXI4DMAO11Ol
,
CAXI4DMAI11Ol
,
CAXI4DMAOIOOI
,
CAXI4DMAl11Ol
,
CAXI4DMAOOOIl
,
CAXI4DMAllllI
,
CAXI4DMAII0OI
,
CAXI4DMAlI0OI
,
CAXI4DMAI1IlI
,
CAXI4DMAIOOIl
,
CAXI4DMAlOOIl
,
CAXI4DMAOIOIl
,
CAXI4DMAIIOIl
,
CAXI4DMAlIOIl
,
CAXI4DMAOlOIl
,
CAXI4DMAIlOIl
)
;
parameter
NUM_INT_BDS
=
0
;
parameter
CAXI4DMAOIO1
=
5
;
parameter
NUM_PRI_LVLS
=
1
;
parameter
CAXI4DMAl0OI
=
23
;
input
CAXI4DMAI
;
input
CAXI4DMAl
;
input
CAXI4DMAIlllI
;
input
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI0llI
;
input
CAXI4DMAOIl1I
;
input
[
31
:
0
]
CAXI4DMAlOl1I
;
input
CAXI4DMAIIl1I
;
input
[
31
:
0
]
CAXI4DMAOll1I
;
input
[
1
:
0
]
CAXI4DMAIll1I
;
input
[
2
:
0
]
CAXI4DMAlll1I
;
input
[
2
:
0
]
CAXI4DMAOO01I
;
input
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAO0l1I
;
input
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAl100I
;
input
CAXI4DMAI0l1I
;
input
CAXI4DMAl0l1I
;
input
[
31
:
0
]
CAXI4DMAO1l1I
;
input
CAXI4DMAl01Ol
;
input
[
1
:
0
]
CAXI4DMAl1OOl
;
input
CAXI4DMAl1l1
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAO11Ol
;
output
reg
[
CAXI4DMAOIO1
-
1
:
0
]
CAXI4DMAI11Ol
;
output
CAXI4DMAOIOOI
;
output
CAXI4DMAl11Ol
;
output
CAXI4DMAOOOIl
;
output
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAllllI
;
output
CAXI4DMAII0OI
;
output
[
31
:
0
]
CAXI4DMAlI0OI
;
output
CAXI4DMAI1IlI
;
output
[
1
:
0
]
CAXI4DMAIOOIl
;
output
[
2
:
0
]
CAXI4DMAlOOIl
;
output
[
2
:
0
]
CAXI4DMAOIOIl
;
output
[
31
:
0
]
CAXI4DMAIIOIl
;
output
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAlIOIl
;
output
CAXI4DMAOlOIl
;
output
[
31
:
0
]
CAXI4DMAIlOIl
;
reg
[
1
:
0
]
CAXI4DMAIO10l
;
reg
CAXI4DMAlO10l
;
reg
[
31
:
0
]
CAXI4DMAOI10l
;
reg
CAXI4DMAII10l
;
reg
[
31
:
0
]
CAXI4DMAlI10l
;
reg
[
1
:
0
]
CAXI4DMAOl10l
;
reg
[
2
:
0
]
CAXI4DMAIl10l
;
reg
[
2
:
0
]
CAXI4DMAll10l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAO010l
;
reg
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAI010l
;
reg
CAXI4DMAl010l
;
reg
CAXI4DMAO110l
;
reg
[
31
:
0
]
CAXI4DMAI110l
;
reg
CAXI4DMAl110l
;
reg
[
31
:
0
]
CAXI4DMAOOO1l
;
reg
CAXI4DMAIOO1l
;
reg
[
31
:
0
]
CAXI4DMAlOO1l
;
reg
[
1
:
0
]
CAXI4DMAOIO1l
;
reg
[
2
:
0
]
CAXI4DMAIIO1l
;
reg
[
2
:
0
]
CAXI4DMAlIO1l
;
reg
[
CAXI4DMAl0OI
-
1
:
0
]
CAXI4DMAOlO1l
;
reg
[
NUM_PRI_LVLS
-
1
:
0
]
CAXI4DMAIlO1l
;
reg
CAXI4DMAllO1l
;
reg
CAXI4DMAO0O1l
;
reg
[
31
:
0
]
CAXI4DMAI0O1l
;
reg
CAXI4DMAl0O1l
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAIO10l
<=
2
'b
0
;
end
else
begin
case
(
{
CAXI4DMAIlllI
,
CAXI4DMAl1OOl
[
1
]
,
CAXI4DMAl1OOl
[
0
]
}
)
3
'b
000
,
3
'b
101
,
3
'b
110
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
;
end
3
'b
001
,
3
'b
010
,
3
'b
111
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
-
1
'b
1
;
end
3
'b
011
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
-
2
'b
10
;
end
3
'b
100
:
begin
CAXI4DMAIO10l
<=
CAXI4DMAIO10l
+
1
'b
1
;
end
endcase
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAl0O1l
<=
1
'b
0
;
end
else
if
(
CAXI4DMAIlllI
)
begin
CAXI4DMAl0O1l
<=
~
CAXI4DMAl0O1l
;
end
end
assign
CAXI4DMAOlOIl
=
(
CAXI4DMAIO10l
<
2
'b
10
)
?
1
'b
1
:
1
'b
0
;
assign
CAXI4DMAOOOIl
=
(
CAXI4DMAIO10l
!=
2
'b
0
)
;
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAO11Ol
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAlO10l
<=
1
'b
0
;
CAXI4DMAOI10l
<=
32
'b
0
;
CAXI4DMAII10l
<=
1
'b
0
;
CAXI4DMAlI10l
<=
32
'b
0
;
CAXI4DMAOl10l
<=
2
'b
0
;
CAXI4DMAIl10l
<=
3
'b
0
;
CAXI4DMAll10l
<=
3
'b
0
;
CAXI4DMAO010l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAI010l
<=
{
NUM_PRI_LVLS
{
1
'b
0
}
}
;
CAXI4DMAl010l
<=
1
'b
0
;
CAXI4DMAO110l
<=
1
'b
0
;
CAXI4DMAI110l
<=
32
'b
0
;
end
else
begin
if
(
CAXI4DMAIlllI
&
!
CAXI4DMAl0O1l
)
begin
CAXI4DMAO11Ol
<=
CAXI4DMAI0llI
;
CAXI4DMAlO10l
<=
CAXI4DMAOIl1I
;
CAXI4DMAOI10l
<=
CAXI4DMAlOl1I
;
CAXI4DMAII10l
<=
CAXI4DMAIIl1I
;
CAXI4DMAlI10l
<=
CAXI4DMAOll1I
;
CAXI4DMAOl10l
<=
CAXI4DMAIll1I
;
CAXI4DMAIl10l
<=
CAXI4DMAlll1I
;
CAXI4DMAll10l
<=
CAXI4DMAOO01I
;
CAXI4DMAO010l
<=
CAXI4DMAO0l1I
;
CAXI4DMAI010l
<=
CAXI4DMAl100I
;
CAXI4DMAl010l
<=
CAXI4DMAI0l1I
;
CAXI4DMAO110l
<=
CAXI4DMAl0l1I
;
CAXI4DMAI110l
<=
CAXI4DMAO1l1I
;
end
end
end
always
@
(
posedge
CAXI4DMAI
or
negedge
CAXI4DMAl
)
begin
if
(
!
CAXI4DMAl
)
begin
CAXI4DMAI11Ol
<=
{
CAXI4DMAOIO1
{
1
'b
0
}
}
;
CAXI4DMAl110l
<=
1
'b
0
;
CAXI4DMAOOO1l
<=
32
'b
0
;
CAXI4DMAIOO1l
<=
1
'b
0
;
CAXI4DMAlOO1l
<=
32
'b
0
;
CAXI4DMAOIO1l
<=
2
'b
0
;
CAXI4DMAIIO1l
<=
3
'b
0
;
CAXI4DMAlIO1l
<=
3
'b
0
;
CAXI4DMAOlO1l
<=
{
CAXI4DMAl0OI
{
1
'b
0
}
}
;
CAXI4DMAIlO1l
<=
{
NUM_PRI_LVLS
{
1
'b
0
}
}
;
CAXI4DMAllO1l
<=
1
'b
0
;
CAXI4DMAO0O1l
<=
1
'b
0
;
CAXI4DMAI0O1l
<=
32
'b
0
;
end
else
begin
if
(
CAXI4DMAIlllI
&
CAXI4DMAl0O1l
)
begin
CAXI4DMAI11Ol
<=
CAXI4DMAI0llI
;
CAXI4DMAl110l
<=
CAXI4DMAOIl1I
;
CAXI4DMAOOO1l
<=
CAXI4DMAlOl1I
;
CAXI4DMAIOO1l
<=
CAXI4DMAIIl1I
;
CAXI4DMAlOO1l
<=
CAXI4DMAOll1I
;
CAXI4DMAOIO1l
<=
CAXI4DMAIll1I
;
CAXI4DMAIIO1l
<=
CAXI4DMAlll1I
;
CAXI4DMAlIO1l
<=
CAXI4DMAOO01I
;
CAXI4DMAOlO1l
<=
CAXI4DMAO0l1I
;
CAXI4DMAIlO1l
<=
CAXI4DMAl100I
;
CAXI4DMAllO1l
<=
CAXI4DMAI0l1I
;
CAXI4DMAO0O1l
<=
CAXI4DMAl0l1I
;
CAXI4DMAI0O1l
<=
CAXI4DMAO1l1I
;
end
end
end
assign
CAXI4DMAII0OI
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAl110l
:
CAXI4DMAOI10l
;
assign
CAXI4DMAlI0OI
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAOOO1l
:
CAXI4DMAOI10l
;
assign
CAXI4DMAI1IlI
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAIOO1l
:
CAXI4DMAII10l
;
assign
CAXI4DMAIOOIl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAOIO1l
:
CAXI4DMAOl10l
;
assign
CAXI4DMAlOOIl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAIIO1l
:
CAXI4DMAIl10l
;
assign
CAXI4DMAOIOIl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAlIO1l
:
CAXI4DMAll10l
;
assign
CAXI4DMAIIOIl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAlOO1l
:
CAXI4DMAlI10l
;
assign
CAXI4DMAlIOIl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAOlO1l
:
CAXI4DMAO010l
;
assign
CAXI4DMAllllI
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAIlO1l
:
CAXI4DMAI010l
;
assign
CAXI4DMAOIOOI
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAllO1l
:
CAXI4DMAl010l
;
assign
CAXI4DMAl11Ol
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAO0O1l
:
CAXI4DMAO110l
;
assign
CAXI4DMAIlOIl
=
(
CAXI4DMAl1l1
)
?
CAXI4DMAI0O1l
:
CAXI4DMAI110l
;
endmodule
